//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul  7 20:54:34 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_1__0_ -----
module sb_1__0_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:295] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:295] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:295] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:295] chany_top_out;
//----- OUTPUT PORTS -----
output [0:295] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:295] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_33_sram;
wire [0:1] mux_tree_tapbuf_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_34_sram;
wire [0:1] mux_tree_tapbuf_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_35_sram;
wire [0:1] mux_tree_tapbuf_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_36_sram;
wire [0:1] mux_tree_tapbuf_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_37_sram;
wire [0:1] mux_tree_tapbuf_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_38_sram;
wire [0:1] mux_tree_tapbuf_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_39_sram;
wire [0:1] mux_tree_tapbuf_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_40_sram;
wire [0:1] mux_tree_tapbuf_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_41_sram;
wire [0:1] mux_tree_tapbuf_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_42_sram;
wire [0:1] mux_tree_tapbuf_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_43_sram;
wire [0:1] mux_tree_tapbuf_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_44_sram;
wire [0:1] mux_tree_tapbuf_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_45_sram;
wire [0:1] mux_tree_tapbuf_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_46_sram;
wire [0:1] mux_tree_tapbuf_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_47_sram;
wire [0:1] mux_tree_tapbuf_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_48_sram;
wire [0:1] mux_tree_tapbuf_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_49_sram;
wire [0:1] mux_tree_tapbuf_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_50_sram;
wire [0:1] mux_tree_tapbuf_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_51_sram;
wire [0:1] mux_tree_tapbuf_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_52_sram;
wire [0:1] mux_tree_tapbuf_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_53_sram;
wire [0:1] mux_tree_tapbuf_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_54_sram;
wire [0:1] mux_tree_tapbuf_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_55_sram;
wire [0:1] mux_tree_tapbuf_size3_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_56_sram;
wire [0:1] mux_tree_tapbuf_size3_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_57_sram;
wire [0:1] mux_tree_tapbuf_size3_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_58_sram;
wire [0:1] mux_tree_tapbuf_size3_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_59_sram;
wire [0:1] mux_tree_tapbuf_size3_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_60_sram;
wire [0:1] mux_tree_tapbuf_size3_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_61_sram;
wire [0:1] mux_tree_tapbuf_size3_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_62_sram;
wire [0:1] mux_tree_tapbuf_size3_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_63_sram;
wire [0:1] mux_tree_tapbuf_size3_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_64_sram;
wire [0:1] mux_tree_tapbuf_size3_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_65_sram;
wire [0:1] mux_tree_tapbuf_size3_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_66_sram;
wire [0:1] mux_tree_tapbuf_size3_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_100_sram;
wire [0:2] mux_tree_tapbuf_size4_100_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_101_sram;
wire [0:2] mux_tree_tapbuf_size4_101_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_102_sram;
wire [0:2] mux_tree_tapbuf_size4_102_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_103_sram;
wire [0:2] mux_tree_tapbuf_size4_103_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_104_sram;
wire [0:2] mux_tree_tapbuf_size4_104_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_105_sram;
wire [0:2] mux_tree_tapbuf_size4_105_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_106_sram;
wire [0:2] mux_tree_tapbuf_size4_106_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_107_sram;
wire [0:2] mux_tree_tapbuf_size4_107_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_108_sram;
wire [0:2] mux_tree_tapbuf_size4_108_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_109_sram;
wire [0:2] mux_tree_tapbuf_size4_109_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_10_sram;
wire [0:2] mux_tree_tapbuf_size4_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_110_sram;
wire [0:2] mux_tree_tapbuf_size4_110_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_111_sram;
wire [0:2] mux_tree_tapbuf_size4_111_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_112_sram;
wire [0:2] mux_tree_tapbuf_size4_112_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_113_sram;
wire [0:2] mux_tree_tapbuf_size4_113_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_114_sram;
wire [0:2] mux_tree_tapbuf_size4_114_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_115_sram;
wire [0:2] mux_tree_tapbuf_size4_115_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_116_sram;
wire [0:2] mux_tree_tapbuf_size4_116_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_117_sram;
wire [0:2] mux_tree_tapbuf_size4_117_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_118_sram;
wire [0:2] mux_tree_tapbuf_size4_118_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_119_sram;
wire [0:2] mux_tree_tapbuf_size4_119_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_11_sram;
wire [0:2] mux_tree_tapbuf_size4_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_120_sram;
wire [0:2] mux_tree_tapbuf_size4_120_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_121_sram;
wire [0:2] mux_tree_tapbuf_size4_121_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_122_sram;
wire [0:2] mux_tree_tapbuf_size4_122_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_123_sram;
wire [0:2] mux_tree_tapbuf_size4_123_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_124_sram;
wire [0:2] mux_tree_tapbuf_size4_124_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_125_sram;
wire [0:2] mux_tree_tapbuf_size4_125_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_126_sram;
wire [0:2] mux_tree_tapbuf_size4_126_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_127_sram;
wire [0:2] mux_tree_tapbuf_size4_127_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_128_sram;
wire [0:2] mux_tree_tapbuf_size4_128_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_129_sram;
wire [0:2] mux_tree_tapbuf_size4_129_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_12_sram;
wire [0:2] mux_tree_tapbuf_size4_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_130_sram;
wire [0:2] mux_tree_tapbuf_size4_130_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_131_sram;
wire [0:2] mux_tree_tapbuf_size4_131_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_132_sram;
wire [0:2] mux_tree_tapbuf_size4_132_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_133_sram;
wire [0:2] mux_tree_tapbuf_size4_133_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_134_sram;
wire [0:2] mux_tree_tapbuf_size4_134_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_135_sram;
wire [0:2] mux_tree_tapbuf_size4_135_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_136_sram;
wire [0:2] mux_tree_tapbuf_size4_136_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_137_sram;
wire [0:2] mux_tree_tapbuf_size4_137_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_138_sram;
wire [0:2] mux_tree_tapbuf_size4_138_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_139_sram;
wire [0:2] mux_tree_tapbuf_size4_139_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_13_sram;
wire [0:2] mux_tree_tapbuf_size4_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_140_sram;
wire [0:2] mux_tree_tapbuf_size4_140_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_141_sram;
wire [0:2] mux_tree_tapbuf_size4_141_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_142_sram;
wire [0:2] mux_tree_tapbuf_size4_142_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_143_sram;
wire [0:2] mux_tree_tapbuf_size4_143_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_144_sram;
wire [0:2] mux_tree_tapbuf_size4_144_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_145_sram;
wire [0:2] mux_tree_tapbuf_size4_145_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_146_sram;
wire [0:2] mux_tree_tapbuf_size4_146_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_147_sram;
wire [0:2] mux_tree_tapbuf_size4_147_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_148_sram;
wire [0:2] mux_tree_tapbuf_size4_148_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_149_sram;
wire [0:2] mux_tree_tapbuf_size4_149_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_14_sram;
wire [0:2] mux_tree_tapbuf_size4_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_150_sram;
wire [0:2] mux_tree_tapbuf_size4_150_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_151_sram;
wire [0:2] mux_tree_tapbuf_size4_151_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_152_sram;
wire [0:2] mux_tree_tapbuf_size4_152_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_153_sram;
wire [0:2] mux_tree_tapbuf_size4_153_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_154_sram;
wire [0:2] mux_tree_tapbuf_size4_154_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_155_sram;
wire [0:2] mux_tree_tapbuf_size4_155_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_156_sram;
wire [0:2] mux_tree_tapbuf_size4_156_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_157_sram;
wire [0:2] mux_tree_tapbuf_size4_157_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_158_sram;
wire [0:2] mux_tree_tapbuf_size4_158_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_159_sram;
wire [0:2] mux_tree_tapbuf_size4_159_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_15_sram;
wire [0:2] mux_tree_tapbuf_size4_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_160_sram;
wire [0:2] mux_tree_tapbuf_size4_160_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_161_sram;
wire [0:2] mux_tree_tapbuf_size4_161_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_162_sram;
wire [0:2] mux_tree_tapbuf_size4_162_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_163_sram;
wire [0:2] mux_tree_tapbuf_size4_163_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_164_sram;
wire [0:2] mux_tree_tapbuf_size4_164_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_165_sram;
wire [0:2] mux_tree_tapbuf_size4_165_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_166_sram;
wire [0:2] mux_tree_tapbuf_size4_166_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_167_sram;
wire [0:2] mux_tree_tapbuf_size4_167_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_168_sram;
wire [0:2] mux_tree_tapbuf_size4_168_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_169_sram;
wire [0:2] mux_tree_tapbuf_size4_169_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_16_sram;
wire [0:2] mux_tree_tapbuf_size4_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_170_sram;
wire [0:2] mux_tree_tapbuf_size4_170_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_171_sram;
wire [0:2] mux_tree_tapbuf_size4_171_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_172_sram;
wire [0:2] mux_tree_tapbuf_size4_172_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_173_sram;
wire [0:2] mux_tree_tapbuf_size4_173_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_174_sram;
wire [0:2] mux_tree_tapbuf_size4_174_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_175_sram;
wire [0:2] mux_tree_tapbuf_size4_175_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_176_sram;
wire [0:2] mux_tree_tapbuf_size4_176_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_177_sram;
wire [0:2] mux_tree_tapbuf_size4_177_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_178_sram;
wire [0:2] mux_tree_tapbuf_size4_178_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_179_sram;
wire [0:2] mux_tree_tapbuf_size4_179_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_17_sram;
wire [0:2] mux_tree_tapbuf_size4_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_180_sram;
wire [0:2] mux_tree_tapbuf_size4_180_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_181_sram;
wire [0:2] mux_tree_tapbuf_size4_181_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_182_sram;
wire [0:2] mux_tree_tapbuf_size4_182_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_183_sram;
wire [0:2] mux_tree_tapbuf_size4_183_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_184_sram;
wire [0:2] mux_tree_tapbuf_size4_184_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_185_sram;
wire [0:2] mux_tree_tapbuf_size4_185_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_186_sram;
wire [0:2] mux_tree_tapbuf_size4_186_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_187_sram;
wire [0:2] mux_tree_tapbuf_size4_187_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_188_sram;
wire [0:2] mux_tree_tapbuf_size4_188_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_189_sram;
wire [0:2] mux_tree_tapbuf_size4_189_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_18_sram;
wire [0:2] mux_tree_tapbuf_size4_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_190_sram;
wire [0:2] mux_tree_tapbuf_size4_190_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_191_sram;
wire [0:2] mux_tree_tapbuf_size4_191_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_192_sram;
wire [0:2] mux_tree_tapbuf_size4_192_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_193_sram;
wire [0:2] mux_tree_tapbuf_size4_193_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_194_sram;
wire [0:2] mux_tree_tapbuf_size4_194_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_195_sram;
wire [0:2] mux_tree_tapbuf_size4_195_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_196_sram;
wire [0:2] mux_tree_tapbuf_size4_196_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_197_sram;
wire [0:2] mux_tree_tapbuf_size4_197_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_198_sram;
wire [0:2] mux_tree_tapbuf_size4_198_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_199_sram;
wire [0:2] mux_tree_tapbuf_size4_199_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_19_sram;
wire [0:2] mux_tree_tapbuf_size4_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_200_sram;
wire [0:2] mux_tree_tapbuf_size4_200_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_201_sram;
wire [0:2] mux_tree_tapbuf_size4_201_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_202_sram;
wire [0:2] mux_tree_tapbuf_size4_202_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_203_sram;
wire [0:2] mux_tree_tapbuf_size4_203_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_204_sram;
wire [0:2] mux_tree_tapbuf_size4_204_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_205_sram;
wire [0:2] mux_tree_tapbuf_size4_205_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_206_sram;
wire [0:2] mux_tree_tapbuf_size4_206_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_207_sram;
wire [0:2] mux_tree_tapbuf_size4_207_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_208_sram;
wire [0:2] mux_tree_tapbuf_size4_208_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_209_sram;
wire [0:2] mux_tree_tapbuf_size4_209_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_20_sram;
wire [0:2] mux_tree_tapbuf_size4_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_210_sram;
wire [0:2] mux_tree_tapbuf_size4_210_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_211_sram;
wire [0:2] mux_tree_tapbuf_size4_211_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_212_sram;
wire [0:2] mux_tree_tapbuf_size4_212_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_213_sram;
wire [0:2] mux_tree_tapbuf_size4_213_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_214_sram;
wire [0:2] mux_tree_tapbuf_size4_214_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_215_sram;
wire [0:2] mux_tree_tapbuf_size4_215_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_216_sram;
wire [0:2] mux_tree_tapbuf_size4_216_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_217_sram;
wire [0:2] mux_tree_tapbuf_size4_217_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_218_sram;
wire [0:2] mux_tree_tapbuf_size4_218_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_219_sram;
wire [0:2] mux_tree_tapbuf_size4_219_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_21_sram;
wire [0:2] mux_tree_tapbuf_size4_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_220_sram;
wire [0:2] mux_tree_tapbuf_size4_220_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_221_sram;
wire [0:2] mux_tree_tapbuf_size4_221_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_222_sram;
wire [0:2] mux_tree_tapbuf_size4_222_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_223_sram;
wire [0:2] mux_tree_tapbuf_size4_223_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_224_sram;
wire [0:2] mux_tree_tapbuf_size4_224_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_225_sram;
wire [0:2] mux_tree_tapbuf_size4_225_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_226_sram;
wire [0:2] mux_tree_tapbuf_size4_226_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_22_sram;
wire [0:2] mux_tree_tapbuf_size4_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_23_sram;
wire [0:2] mux_tree_tapbuf_size4_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_24_sram;
wire [0:2] mux_tree_tapbuf_size4_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_25_sram;
wire [0:2] mux_tree_tapbuf_size4_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_26_sram;
wire [0:2] mux_tree_tapbuf_size4_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_27_sram;
wire [0:2] mux_tree_tapbuf_size4_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_28_sram;
wire [0:2] mux_tree_tapbuf_size4_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_29_sram;
wire [0:2] mux_tree_tapbuf_size4_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_30_sram;
wire [0:2] mux_tree_tapbuf_size4_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_31_sram;
wire [0:2] mux_tree_tapbuf_size4_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_32_sram;
wire [0:2] mux_tree_tapbuf_size4_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_33_sram;
wire [0:2] mux_tree_tapbuf_size4_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_34_sram;
wire [0:2] mux_tree_tapbuf_size4_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_35_sram;
wire [0:2] mux_tree_tapbuf_size4_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_36_sram;
wire [0:2] mux_tree_tapbuf_size4_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_37_sram;
wire [0:2] mux_tree_tapbuf_size4_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_38_sram;
wire [0:2] mux_tree_tapbuf_size4_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_39_sram;
wire [0:2] mux_tree_tapbuf_size4_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_40_sram;
wire [0:2] mux_tree_tapbuf_size4_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_41_sram;
wire [0:2] mux_tree_tapbuf_size4_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_42_sram;
wire [0:2] mux_tree_tapbuf_size4_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_43_sram;
wire [0:2] mux_tree_tapbuf_size4_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_44_sram;
wire [0:2] mux_tree_tapbuf_size4_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_45_sram;
wire [0:2] mux_tree_tapbuf_size4_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_46_sram;
wire [0:2] mux_tree_tapbuf_size4_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_47_sram;
wire [0:2] mux_tree_tapbuf_size4_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_48_sram;
wire [0:2] mux_tree_tapbuf_size4_48_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_49_sram;
wire [0:2] mux_tree_tapbuf_size4_49_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_4_sram;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_50_sram;
wire [0:2] mux_tree_tapbuf_size4_50_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_51_sram;
wire [0:2] mux_tree_tapbuf_size4_51_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_52_sram;
wire [0:2] mux_tree_tapbuf_size4_52_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_53_sram;
wire [0:2] mux_tree_tapbuf_size4_53_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_54_sram;
wire [0:2] mux_tree_tapbuf_size4_54_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_55_sram;
wire [0:2] mux_tree_tapbuf_size4_55_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_56_sram;
wire [0:2] mux_tree_tapbuf_size4_56_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_57_sram;
wire [0:2] mux_tree_tapbuf_size4_57_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_58_sram;
wire [0:2] mux_tree_tapbuf_size4_58_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_59_sram;
wire [0:2] mux_tree_tapbuf_size4_59_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_5_sram;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_60_sram;
wire [0:2] mux_tree_tapbuf_size4_60_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_61_sram;
wire [0:2] mux_tree_tapbuf_size4_61_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_62_sram;
wire [0:2] mux_tree_tapbuf_size4_62_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_63_sram;
wire [0:2] mux_tree_tapbuf_size4_63_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_64_sram;
wire [0:2] mux_tree_tapbuf_size4_64_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_65_sram;
wire [0:2] mux_tree_tapbuf_size4_65_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_66_sram;
wire [0:2] mux_tree_tapbuf_size4_66_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_67_sram;
wire [0:2] mux_tree_tapbuf_size4_67_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_68_sram;
wire [0:2] mux_tree_tapbuf_size4_68_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_69_sram;
wire [0:2] mux_tree_tapbuf_size4_69_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_6_sram;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_70_sram;
wire [0:2] mux_tree_tapbuf_size4_70_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_71_sram;
wire [0:2] mux_tree_tapbuf_size4_71_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_72_sram;
wire [0:2] mux_tree_tapbuf_size4_72_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_73_sram;
wire [0:2] mux_tree_tapbuf_size4_73_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_74_sram;
wire [0:2] mux_tree_tapbuf_size4_74_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_75_sram;
wire [0:2] mux_tree_tapbuf_size4_75_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_76_sram;
wire [0:2] mux_tree_tapbuf_size4_76_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_77_sram;
wire [0:2] mux_tree_tapbuf_size4_77_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_78_sram;
wire [0:2] mux_tree_tapbuf_size4_78_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_79_sram;
wire [0:2] mux_tree_tapbuf_size4_79_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_7_sram;
wire [0:2] mux_tree_tapbuf_size4_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_80_sram;
wire [0:2] mux_tree_tapbuf_size4_80_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_81_sram;
wire [0:2] mux_tree_tapbuf_size4_81_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_82_sram;
wire [0:2] mux_tree_tapbuf_size4_82_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_83_sram;
wire [0:2] mux_tree_tapbuf_size4_83_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_84_sram;
wire [0:2] mux_tree_tapbuf_size4_84_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_85_sram;
wire [0:2] mux_tree_tapbuf_size4_85_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_86_sram;
wire [0:2] mux_tree_tapbuf_size4_86_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_87_sram;
wire [0:2] mux_tree_tapbuf_size4_87_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_88_sram;
wire [0:2] mux_tree_tapbuf_size4_88_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_89_sram;
wire [0:2] mux_tree_tapbuf_size4_89_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_8_sram;
wire [0:2] mux_tree_tapbuf_size4_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_90_sram;
wire [0:2] mux_tree_tapbuf_size4_90_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_91_sram;
wire [0:2] mux_tree_tapbuf_size4_91_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_92_sram;
wire [0:2] mux_tree_tapbuf_size4_92_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_93_sram;
wire [0:2] mux_tree_tapbuf_size4_93_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_94_sram;
wire [0:2] mux_tree_tapbuf_size4_94_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_95_sram;
wire [0:2] mux_tree_tapbuf_size4_95_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_96_sram;
wire [0:2] mux_tree_tapbuf_size4_96_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_97_sram;
wire [0:2] mux_tree_tapbuf_size4_97_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_98_sram;
wire [0:2] mux_tree_tapbuf_size4_98_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_99_sram;
wire [0:2] mux_tree_tapbuf_size4_99_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_9_sram;
wire [0:2] mux_tree_tapbuf_size4_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_136_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_137_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_138_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_139_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_140_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_141_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_142_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_143_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_144_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_145_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_146_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_147_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_148_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_149_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_150_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_151_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_152_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_153_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_154_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_155_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_156_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_157_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_158_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_159_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_160_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_161_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_162_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_163_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_164_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_165_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_166_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_167_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_168_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_169_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_170_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_171_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_172_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_173_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_174_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_175_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_176_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_177_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_178_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_179_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_180_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_181_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_182_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_183_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_184_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_185_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_186_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_187_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_188_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_189_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_190_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_191_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_192_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_193_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_194_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_195_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_196_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_197_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_198_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_199_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_200_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_201_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_202_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_203_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_204_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_205_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_206_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_207_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_208_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_209_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_210_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_211_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_212_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_213_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_214_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_215_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_216_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_217_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_218_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_219_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_220_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_221_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_222_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_223_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_224_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_225_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_226_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_100_sram;
wire [0:2] mux_tree_tapbuf_size6_100_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_10_sram;
wire [0:2] mux_tree_tapbuf_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_11_sram;
wire [0:2] mux_tree_tapbuf_size6_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_12_sram;
wire [0:2] mux_tree_tapbuf_size6_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_13_sram;
wire [0:2] mux_tree_tapbuf_size6_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_14_sram;
wire [0:2] mux_tree_tapbuf_size6_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_15_sram;
wire [0:2] mux_tree_tapbuf_size6_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_16_sram;
wire [0:2] mux_tree_tapbuf_size6_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_17_sram;
wire [0:2] mux_tree_tapbuf_size6_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_18_sram;
wire [0:2] mux_tree_tapbuf_size6_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_19_sram;
wire [0:2] mux_tree_tapbuf_size6_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_20_sram;
wire [0:2] mux_tree_tapbuf_size6_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_21_sram;
wire [0:2] mux_tree_tapbuf_size6_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_22_sram;
wire [0:2] mux_tree_tapbuf_size6_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_23_sram;
wire [0:2] mux_tree_tapbuf_size6_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_24_sram;
wire [0:2] mux_tree_tapbuf_size6_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_25_sram;
wire [0:2] mux_tree_tapbuf_size6_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_26_sram;
wire [0:2] mux_tree_tapbuf_size6_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_27_sram;
wire [0:2] mux_tree_tapbuf_size6_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_28_sram;
wire [0:2] mux_tree_tapbuf_size6_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_29_sram;
wire [0:2] mux_tree_tapbuf_size6_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_30_sram;
wire [0:2] mux_tree_tapbuf_size6_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_31_sram;
wire [0:2] mux_tree_tapbuf_size6_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_32_sram;
wire [0:2] mux_tree_tapbuf_size6_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_33_sram;
wire [0:2] mux_tree_tapbuf_size6_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_34_sram;
wire [0:2] mux_tree_tapbuf_size6_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_35_sram;
wire [0:2] mux_tree_tapbuf_size6_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_36_sram;
wire [0:2] mux_tree_tapbuf_size6_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_37_sram;
wire [0:2] mux_tree_tapbuf_size6_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_38_sram;
wire [0:2] mux_tree_tapbuf_size6_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_39_sram;
wire [0:2] mux_tree_tapbuf_size6_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_40_sram;
wire [0:2] mux_tree_tapbuf_size6_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_41_sram;
wire [0:2] mux_tree_tapbuf_size6_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_42_sram;
wire [0:2] mux_tree_tapbuf_size6_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_43_sram;
wire [0:2] mux_tree_tapbuf_size6_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_44_sram;
wire [0:2] mux_tree_tapbuf_size6_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_45_sram;
wire [0:2] mux_tree_tapbuf_size6_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_46_sram;
wire [0:2] mux_tree_tapbuf_size6_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_47_sram;
wire [0:2] mux_tree_tapbuf_size6_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_48_sram;
wire [0:2] mux_tree_tapbuf_size6_48_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_49_sram;
wire [0:2] mux_tree_tapbuf_size6_49_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_50_sram;
wire [0:2] mux_tree_tapbuf_size6_50_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_51_sram;
wire [0:2] mux_tree_tapbuf_size6_51_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_52_sram;
wire [0:2] mux_tree_tapbuf_size6_52_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_53_sram;
wire [0:2] mux_tree_tapbuf_size6_53_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_54_sram;
wire [0:2] mux_tree_tapbuf_size6_54_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_55_sram;
wire [0:2] mux_tree_tapbuf_size6_55_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_56_sram;
wire [0:2] mux_tree_tapbuf_size6_56_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_57_sram;
wire [0:2] mux_tree_tapbuf_size6_57_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_58_sram;
wire [0:2] mux_tree_tapbuf_size6_58_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_59_sram;
wire [0:2] mux_tree_tapbuf_size6_59_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_60_sram;
wire [0:2] mux_tree_tapbuf_size6_60_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_61_sram;
wire [0:2] mux_tree_tapbuf_size6_61_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_62_sram;
wire [0:2] mux_tree_tapbuf_size6_62_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_63_sram;
wire [0:2] mux_tree_tapbuf_size6_63_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_64_sram;
wire [0:2] mux_tree_tapbuf_size6_64_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_65_sram;
wire [0:2] mux_tree_tapbuf_size6_65_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_66_sram;
wire [0:2] mux_tree_tapbuf_size6_66_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_67_sram;
wire [0:2] mux_tree_tapbuf_size6_67_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_68_sram;
wire [0:2] mux_tree_tapbuf_size6_68_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_69_sram;
wire [0:2] mux_tree_tapbuf_size6_69_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_70_sram;
wire [0:2] mux_tree_tapbuf_size6_70_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_71_sram;
wire [0:2] mux_tree_tapbuf_size6_71_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_72_sram;
wire [0:2] mux_tree_tapbuf_size6_72_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_73_sram;
wire [0:2] mux_tree_tapbuf_size6_73_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_74_sram;
wire [0:2] mux_tree_tapbuf_size6_74_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_75_sram;
wire [0:2] mux_tree_tapbuf_size6_75_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_76_sram;
wire [0:2] mux_tree_tapbuf_size6_76_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_77_sram;
wire [0:2] mux_tree_tapbuf_size6_77_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_78_sram;
wire [0:2] mux_tree_tapbuf_size6_78_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_79_sram;
wire [0:2] mux_tree_tapbuf_size6_79_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_80_sram;
wire [0:2] mux_tree_tapbuf_size6_80_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_81_sram;
wire [0:2] mux_tree_tapbuf_size6_81_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_82_sram;
wire [0:2] mux_tree_tapbuf_size6_82_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_83_sram;
wire [0:2] mux_tree_tapbuf_size6_83_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_84_sram;
wire [0:2] mux_tree_tapbuf_size6_84_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_85_sram;
wire [0:2] mux_tree_tapbuf_size6_85_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_86_sram;
wire [0:2] mux_tree_tapbuf_size6_86_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_87_sram;
wire [0:2] mux_tree_tapbuf_size6_87_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_88_sram;
wire [0:2] mux_tree_tapbuf_size6_88_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_89_sram;
wire [0:2] mux_tree_tapbuf_size6_89_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_90_sram;
wire [0:2] mux_tree_tapbuf_size6_90_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_91_sram;
wire [0:2] mux_tree_tapbuf_size6_91_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_92_sram;
wire [0:2] mux_tree_tapbuf_size6_92_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_93_sram;
wire [0:2] mux_tree_tapbuf_size6_93_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_94_sram;
wire [0:2] mux_tree_tapbuf_size6_94_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_95_sram;
wire [0:2] mux_tree_tapbuf_size6_95_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_96_sram;
wire [0:2] mux_tree_tapbuf_size6_96_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_97_sram;
wire [0:2] mux_tree_tapbuf_size6_97_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_98_sram;
wire [0:2] mux_tree_tapbuf_size6_98_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_99_sram;
wire [0:2] mux_tree_tapbuf_size6_99_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_9_sram;
wire [0:2] mux_tree_tapbuf_size6_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_10_sram;
wire [0:2] mux_tree_tapbuf_size7_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_11_sram;
wire [0:2] mux_tree_tapbuf_size7_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_12_sram;
wire [0:2] mux_tree_tapbuf_size7_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_13_sram;
wire [0:2] mux_tree_tapbuf_size7_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_14_sram;
wire [0:2] mux_tree_tapbuf_size7_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_15_sram;
wire [0:2] mux_tree_tapbuf_size7_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_16_sram;
wire [0:2] mux_tree_tapbuf_size7_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_17_sram;
wire [0:2] mux_tree_tapbuf_size7_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_18_sram;
wire [0:2] mux_tree_tapbuf_size7_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_19_sram;
wire [0:2] mux_tree_tapbuf_size7_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_3_sram;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_4_sram;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_5_sram;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_6_sram;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_7_sram;
wire [0:2] mux_tree_tapbuf_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_8_sram;
wire [0:2] mux_tree_tapbuf_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_9_sram;
wire [0:2] mux_tree_tapbuf_size7_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[150] = chanx_right_in[149];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[151] = chanx_right_in[150];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[153] = chanx_right_in[152];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[154] = chanx_right_in[153];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[155] = chanx_right_in[154];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[157] = chanx_right_in[156];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[158] = chanx_right_in[157];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[159] = chanx_right_in[158];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[161] = chanx_right_in[160];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[162] = chanx_right_in[161];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[163] = chanx_right_in[162];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[165] = chanx_right_in[164];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[166] = chanx_right_in[165];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[167] = chanx_right_in[166];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[169] = chanx_right_in[168];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[170] = chanx_right_in[169];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[171] = chanx_right_in[170];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[173] = chanx_right_in[172];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[174] = chanx_right_in[173];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[175] = chanx_right_in[174];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[177] = chanx_right_in[176];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[178] = chanx_right_in[177];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[179] = chanx_right_in[178];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[181] = chanx_right_in[180];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[182] = chanx_right_in[181];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[183] = chanx_right_in[182];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[185] = chanx_right_in[184];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[186] = chanx_right_in[185];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[187] = chanx_right_in[186];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[189] = chanx_right_in[188];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[190] = chanx_right_in[189];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[191] = chanx_right_in[190];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[193] = chanx_right_in[192];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[194] = chanx_right_in[193];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[195] = chanx_right_in[194];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[197] = chanx_right_in[196];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[198] = chanx_right_in[197];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[199] = chanx_right_in[198];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[201] = chanx_right_in[200];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[202] = chanx_right_in[201];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[203] = chanx_right_in[202];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[205] = chanx_right_in[204];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[206] = chanx_right_in[205];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[207] = chanx_right_in[206];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[209] = chanx_right_in[208];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[210] = chanx_right_in[209];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[211] = chanx_right_in[210];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[213] = chanx_right_in[212];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[214] = chanx_right_in[213];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[215] = chanx_right_in[214];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[217] = chanx_right_in[216];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[218] = chanx_right_in[217];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[219] = chanx_right_in[218];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[221] = chanx_right_in[220];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[222] = chanx_right_in[221];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[223] = chanx_right_in[222];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[225] = chanx_right_in[224];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[226] = chanx_right_in[225];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[227] = chanx_right_in[226];
// ----- Local connection due to Wire 540 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[229] = chanx_right_in[228];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[230] = chanx_right_in[229];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[231] = chanx_right_in[230];
// ----- Local connection due to Wire 544 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[233] = chanx_right_in[232];
// ----- Local connection due to Wire 545 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[234] = chanx_right_in[233];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[235] = chanx_right_in[234];
// ----- Local connection due to Wire 548 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[237] = chanx_right_in[236];
// ----- Local connection due to Wire 549 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[238] = chanx_right_in[237];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[239] = chanx_right_in[238];
// ----- Local connection due to Wire 552 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[241] = chanx_right_in[240];
// ----- Local connection due to Wire 553 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[242] = chanx_right_in[241];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[243] = chanx_right_in[242];
// ----- Local connection due to Wire 556 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[245] = chanx_right_in[244];
// ----- Local connection due to Wire 557 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[246] = chanx_right_in[245];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[247] = chanx_right_in[246];
// ----- Local connection due to Wire 560 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[249] = chanx_right_in[248];
// ----- Local connection due to Wire 561 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[250] = chanx_right_in[249];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[251] = chanx_right_in[250];
// ----- Local connection due to Wire 564 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[253] = chanx_right_in[252];
// ----- Local connection due to Wire 565 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[254] = chanx_right_in[253];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[255] = chanx_right_in[254];
// ----- Local connection due to Wire 568 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[257] = chanx_right_in[256];
// ----- Local connection due to Wire 569 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[258] = chanx_right_in[257];
// ----- Local connection due to Wire 570 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[259] = chanx_right_in[258];
// ----- Local connection due to Wire 572 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[261] = chanx_right_in[260];
// ----- Local connection due to Wire 573 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[262] = chanx_right_in[261];
// ----- Local connection due to Wire 574 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[263] = chanx_right_in[262];
// ----- Local connection due to Wire 576 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[265] = chanx_right_in[264];
// ----- Local connection due to Wire 577 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[266] = chanx_right_in[265];
// ----- Local connection due to Wire 578 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[267] = chanx_right_in[266];
// ----- Local connection due to Wire 580 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[269] = chanx_right_in[268];
// ----- Local connection due to Wire 581 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[270] = chanx_right_in[269];
// ----- Local connection due to Wire 582 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[271] = chanx_right_in[270];
// ----- Local connection due to Wire 584 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[273] = chanx_right_in[272];
// ----- Local connection due to Wire 585 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[274] = chanx_right_in[273];
// ----- Local connection due to Wire 586 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[275] = chanx_right_in[274];
// ----- Local connection due to Wire 588 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[277] = chanx_right_in[276];
// ----- Local connection due to Wire 589 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[278] = chanx_right_in[277];
// ----- Local connection due to Wire 590 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[279] = chanx_right_in[278];
// ----- Local connection due to Wire 592 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[281] = chanx_right_in[280];
// ----- Local connection due to Wire 593 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[282] = chanx_right_in[281];
// ----- Local connection due to Wire 594 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[283] = chanx_right_in[282];
// ----- Local connection due to Wire 596 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[285] = chanx_right_in[284];
// ----- Local connection due to Wire 597 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[286] = chanx_right_in[285];
// ----- Local connection due to Wire 598 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[287] = chanx_right_in[286];
// ----- Local connection due to Wire 600 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[289] = chanx_right_in[288];
// ----- Local connection due to Wire 601 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[290] = chanx_right_in[289];
// ----- Local connection due to Wire 602 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[291] = chanx_right_in[290];
// ----- Local connection due to Wire 604 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[293] = chanx_right_in[292];
// ----- Local connection due to Wire 605 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[294] = chanx_right_in[293];
// ----- Local connection due to Wire 606 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[295] = chanx_right_in[294];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 625 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 673 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 674 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 677 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 678 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 681 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 682 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 685 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 686 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 689 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 690 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 693 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 694 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 697 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 698 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 701 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 702 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 705 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 706 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 709 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 710 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 712 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 713 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 714 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 716 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 717 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 718 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 720 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 721 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 722 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 724 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 725 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 726 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 728 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 729 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 730 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 732 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 733 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 734 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 736 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 737 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 738 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 740 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 741 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 742 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 744 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 745 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 746 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 748 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 749 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 750 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 752 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 753 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 754 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 756 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 757 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 758 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 760 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 761 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 762 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 764 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 765 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 766 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 768 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 769 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 770 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 772 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- Local connection due to Wire 773 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[150] = chanx_left_in[149];
// ----- Local connection due to Wire 774 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[150];
// ----- Local connection due to Wire 776 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[153] = chanx_left_in[152];
// ----- Local connection due to Wire 777 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[154] = chanx_left_in[153];
// ----- Local connection due to Wire 778 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[154];
// ----- Local connection due to Wire 780 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[157] = chanx_left_in[156];
// ----- Local connection due to Wire 781 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[158] = chanx_left_in[157];
// ----- Local connection due to Wire 782 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[158];
// ----- Local connection due to Wire 784 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[161] = chanx_left_in[160];
// ----- Local connection due to Wire 785 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[162] = chanx_left_in[161];
// ----- Local connection due to Wire 786 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[163] = chanx_left_in[162];
// ----- Local connection due to Wire 788 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[165] = chanx_left_in[164];
// ----- Local connection due to Wire 789 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[166] = chanx_left_in[165];
// ----- Local connection due to Wire 790 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[167] = chanx_left_in[166];
// ----- Local connection due to Wire 792 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[169] = chanx_left_in[168];
// ----- Local connection due to Wire 793 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[170] = chanx_left_in[169];
// ----- Local connection due to Wire 794 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[171] = chanx_left_in[170];
// ----- Local connection due to Wire 796 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[173] = chanx_left_in[172];
// ----- Local connection due to Wire 797 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[174] = chanx_left_in[173];
// ----- Local connection due to Wire 798 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[175] = chanx_left_in[174];
// ----- Local connection due to Wire 800 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[177] = chanx_left_in[176];
// ----- Local connection due to Wire 801 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[178] = chanx_left_in[177];
// ----- Local connection due to Wire 802 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[179] = chanx_left_in[178];
// ----- Local connection due to Wire 804 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[181] = chanx_left_in[180];
// ----- Local connection due to Wire 805 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[182] = chanx_left_in[181];
// ----- Local connection due to Wire 806 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[183] = chanx_left_in[182];
// ----- Local connection due to Wire 808 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[185] = chanx_left_in[184];
// ----- Local connection due to Wire 809 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[186] = chanx_left_in[185];
// ----- Local connection due to Wire 810 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[187] = chanx_left_in[186];
// ----- Local connection due to Wire 812 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[189] = chanx_left_in[188];
// ----- Local connection due to Wire 813 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[190] = chanx_left_in[189];
// ----- Local connection due to Wire 814 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[191] = chanx_left_in[190];
// ----- Local connection due to Wire 816 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[193] = chanx_left_in[192];
// ----- Local connection due to Wire 817 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[194] = chanx_left_in[193];
// ----- Local connection due to Wire 818 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[195] = chanx_left_in[194];
// ----- Local connection due to Wire 820 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[197] = chanx_left_in[196];
// ----- Local connection due to Wire 821 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[198] = chanx_left_in[197];
// ----- Local connection due to Wire 822 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[199] = chanx_left_in[198];
// ----- Local connection due to Wire 824 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[201] = chanx_left_in[200];
// ----- Local connection due to Wire 825 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[202] = chanx_left_in[201];
// ----- Local connection due to Wire 826 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[203] = chanx_left_in[202];
// ----- Local connection due to Wire 828 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[205] = chanx_left_in[204];
// ----- Local connection due to Wire 829 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[206] = chanx_left_in[205];
// ----- Local connection due to Wire 830 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[207] = chanx_left_in[206];
// ----- Local connection due to Wire 832 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[209] = chanx_left_in[208];
// ----- Local connection due to Wire 833 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[210] = chanx_left_in[209];
// ----- Local connection due to Wire 834 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[211] = chanx_left_in[210];
// ----- Local connection due to Wire 836 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[213] = chanx_left_in[212];
// ----- Local connection due to Wire 837 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[214] = chanx_left_in[213];
// ----- Local connection due to Wire 838 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[215] = chanx_left_in[214];
// ----- Local connection due to Wire 840 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[217] = chanx_left_in[216];
// ----- Local connection due to Wire 841 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[218] = chanx_left_in[217];
// ----- Local connection due to Wire 842 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[219] = chanx_left_in[218];
// ----- Local connection due to Wire 844 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[221] = chanx_left_in[220];
// ----- Local connection due to Wire 845 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[222] = chanx_left_in[221];
// ----- Local connection due to Wire 846 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[223] = chanx_left_in[222];
// ----- Local connection due to Wire 848 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[225] = chanx_left_in[224];
// ----- Local connection due to Wire 849 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[226] = chanx_left_in[225];
// ----- Local connection due to Wire 850 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[227] = chanx_left_in[226];
// ----- Local connection due to Wire 852 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[229] = chanx_left_in[228];
// ----- Local connection due to Wire 853 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[230] = chanx_left_in[229];
// ----- Local connection due to Wire 854 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[231] = chanx_left_in[230];
// ----- Local connection due to Wire 856 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[233] = chanx_left_in[232];
// ----- Local connection due to Wire 857 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[234] = chanx_left_in[233];
// ----- Local connection due to Wire 858 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[235] = chanx_left_in[234];
// ----- Local connection due to Wire 860 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[237] = chanx_left_in[236];
// ----- Local connection due to Wire 861 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[238] = chanx_left_in[237];
// ----- Local connection due to Wire 862 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[239] = chanx_left_in[238];
// ----- Local connection due to Wire 864 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[241] = chanx_left_in[240];
// ----- Local connection due to Wire 865 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[242] = chanx_left_in[241];
// ----- Local connection due to Wire 866 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[243] = chanx_left_in[242];
// ----- Local connection due to Wire 868 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[245] = chanx_left_in[244];
// ----- Local connection due to Wire 869 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[246] = chanx_left_in[245];
// ----- Local connection due to Wire 870 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[247] = chanx_left_in[246];
// ----- Local connection due to Wire 872 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[249] = chanx_left_in[248];
// ----- Local connection due to Wire 873 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[250] = chanx_left_in[249];
// ----- Local connection due to Wire 874 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[251] = chanx_left_in[250];
// ----- Local connection due to Wire 876 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[253] = chanx_left_in[252];
// ----- Local connection due to Wire 877 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[254] = chanx_left_in[253];
// ----- Local connection due to Wire 878 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[255] = chanx_left_in[254];
// ----- Local connection due to Wire 880 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[257] = chanx_left_in[256];
// ----- Local connection due to Wire 881 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[258] = chanx_left_in[257];
// ----- Local connection due to Wire 882 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[259] = chanx_left_in[258];
// ----- Local connection due to Wire 884 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[261] = chanx_left_in[260];
// ----- Local connection due to Wire 885 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[262] = chanx_left_in[261];
// ----- Local connection due to Wire 886 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[263] = chanx_left_in[262];
// ----- Local connection due to Wire 888 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[265] = chanx_left_in[264];
// ----- Local connection due to Wire 889 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[266] = chanx_left_in[265];
// ----- Local connection due to Wire 890 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[267] = chanx_left_in[266];
// ----- Local connection due to Wire 892 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[269] = chanx_left_in[268];
// ----- Local connection due to Wire 893 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[270] = chanx_left_in[269];
// ----- Local connection due to Wire 894 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[271] = chanx_left_in[270];
// ----- Local connection due to Wire 896 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[273] = chanx_left_in[272];
// ----- Local connection due to Wire 897 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[274] = chanx_left_in[273];
// ----- Local connection due to Wire 898 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[275] = chanx_left_in[274];
// ----- Local connection due to Wire 900 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[277] = chanx_left_in[276];
// ----- Local connection due to Wire 901 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[278] = chanx_left_in[277];
// ----- Local connection due to Wire 902 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[279] = chanx_left_in[278];
// ----- Local connection due to Wire 904 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[281] = chanx_left_in[280];
// ----- Local connection due to Wire 905 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[282] = chanx_left_in[281];
// ----- Local connection due to Wire 906 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[283] = chanx_left_in[282];
// ----- Local connection due to Wire 908 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[285] = chanx_left_in[284];
// ----- Local connection due to Wire 909 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[286] = chanx_left_in[285];
// ----- Local connection due to Wire 910 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[287] = chanx_left_in[286];
// ----- Local connection due to Wire 912 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[289] = chanx_left_in[288];
// ----- Local connection due to Wire 913 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[290] = chanx_left_in[289];
// ----- Local connection due to Wire 914 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[291] = chanx_left_in[290];
// ----- Local connection due to Wire 916 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[293] = chanx_left_in[292];
// ----- Local connection due to Wire 917 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[294] = chanx_left_in[293];
// ----- Local connection due to Wire 918 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[295] = chanx_left_in[294];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size6 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[1], chanx_right_in[7], chanx_left_in[0], chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size6 mux_right_track_40 (
		.in({chany_top_in[4], chany_top_in[78], chany_top_in[152], chany_top_in[226], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size6 mux_right_track_48 (
		.in({chany_top_in[5], chany_top_in[79], chany_top_in[153], chany_top_in[227], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size6 mux_right_track_56 (
		.in({chany_top_in[6], chany_top_in[80], chany_top_in[154], chany_top_in[228], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size6 mux_right_track_64 (
		.in({chany_top_in[7], chany_top_in[81], chany_top_in[155], chany_top_in[229], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size6 mux_right_track_112 (
		.in({chany_top_in[13], chany_top_in[87], chany_top_in[161], chany_top_in[235], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size6 mux_right_track_120 (
		.in({chany_top_in[14], chany_top_in[88], chany_top_in[162], chany_top_in[236], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size6 mux_right_track_144 (
		.in({chany_top_in[17], chany_top_in[91], chany_top_in[165], chany_top_in[239], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size6 mux_right_track_152 (
		.in({chany_top_in[18], chany_top_in[92], chany_top_in[166], chany_top_in[240], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size6 mux_right_track_160 (
		.in({chany_top_in[19], chany_top_in[93], chany_top_in[167], chany_top_in[241], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_9_sram_inv[0:2]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size6 mux_right_track_168 (
		.in({chany_top_in[20], chany_top_in[94], chany_top_in[168], chany_top_in[242], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_10_sram_inv[0:2]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size6 mux_right_track_176 (
		.in({chany_top_in[21], chany_top_in[95], chany_top_in[169], chany_top_in[243], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_11_sram_inv[0:2]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size6 mux_right_track_184 (
		.in({chany_top_in[22], chany_top_in[96], chany_top_in[170], chany_top_in[244], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_12_sram_inv[0:2]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size6 mux_right_track_192 (
		.in({chany_top_in[23], chany_top_in[97], chany_top_in[171], chany_top_in[245], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_13_sram_inv[0:2]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size6 mux_right_track_216 (
		.in({chany_top_in[26], chany_top_in[100], chany_top_in[174], chany_top_in[248], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_14_sram_inv[0:2]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size6 mux_right_track_224 (
		.in({chany_top_in[27], chany_top_in[101], chany_top_in[175], chany_top_in[249], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_15_sram_inv[0:2]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size6 mux_right_track_232 (
		.in({chany_top_in[28], chany_top_in[102], chany_top_in[176], chany_top_in[250], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_16_sram_inv[0:2]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size6 mux_right_track_240 (
		.in({chany_top_in[29], chany_top_in[103], chany_top_in[177], chany_top_in[251], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_17_sram_inv[0:2]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size6 mux_right_track_248 (
		.in({chany_top_in[30], chany_top_in[104], chany_top_in[178], chany_top_in[252], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_18_sram_inv[0:2]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size6 mux_right_track_256 (
		.in({chany_top_in[31], chany_top_in[105], chany_top_in[179], chany_top_in[253], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_19_sram_inv[0:2]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size6 mux_right_track_264 (
		.in({chany_top_in[32], chany_top_in[106], chany_top_in[180], chany_top_in[254], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_20_sram_inv[0:2]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size6 mux_right_track_288 (
		.in({chany_top_in[35], chany_top_in[109], chany_top_in[183], chany_top_in[257], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_21_sram_inv[0:2]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size6 mux_right_track_296 (
		.in({chany_top_in[36], chany_top_in[110], chany_top_in[184], chany_top_in[258], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_22_sram_inv[0:2]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size6 mux_right_track_304 (
		.in({chany_top_in[37], chany_top_in[111], chany_top_in[185], chany_top_in[259], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_23_sram_inv[0:2]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size6 mux_right_track_312 (
		.in({chany_top_in[38], chany_top_in[112], chany_top_in[186], chany_top_in[260], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_24_sram_inv[0:2]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size6 mux_right_track_320 (
		.in({chany_top_in[39], chany_top_in[113], chany_top_in[187], chany_top_in[261], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_25_sram_inv[0:2]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size6 mux_right_track_328 (
		.in({chany_top_in[40], chany_top_in[114], chany_top_in[188], chany_top_in[262], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_26_sram_inv[0:2]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size6 mux_right_track_336 (
		.in({chany_top_in[41], chany_top_in[115], chany_top_in[189], chany_top_in[263], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_27_sram_inv[0:2]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size6 mux_right_track_360 (
		.in({chany_top_in[44], chany_top_in[118], chany_top_in[192], chany_top_in[266], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_28_sram_inv[0:2]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size6 mux_right_track_368 (
		.in({chany_top_in[45], chany_top_in[119], chany_top_in[193], chany_top_in[267], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_29_sram_inv[0:2]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size6 mux_right_track_376 (
		.in({chany_top_in[46], chany_top_in[120], chany_top_in[194], chany_top_in[268], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_30_sram_inv[0:2]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size6 mux_right_track_384 (
		.in({chany_top_in[47], chany_top_in[121], chany_top_in[195], chany_top_in[269], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_31_sram_inv[0:2]),
		.out(chanx_right_out[192]));

	mux_tree_tapbuf_size6 mux_right_track_392 (
		.in({chany_top_in[48], chany_top_in[122], chany_top_in[196], chany_top_in[270], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_32_sram_inv[0:2]),
		.out(chanx_right_out[196]));

	mux_tree_tapbuf_size6 mux_right_track_400 (
		.in({chany_top_in[49], chany_top_in[123], chany_top_in[197], chany_top_in[271], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_33_sram_inv[0:2]),
		.out(chanx_right_out[200]));

	mux_tree_tapbuf_size6 mux_right_track_408 (
		.in({chany_top_in[50], chany_top_in[124], chany_top_in[198], chany_top_in[272], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_34_sram_inv[0:2]),
		.out(chanx_right_out[204]));

	mux_tree_tapbuf_size6 mux_right_track_432 (
		.in({chany_top_in[53], chany_top_in[127], chany_top_in[201], chany_top_in[275], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_35_sram_inv[0:2]),
		.out(chanx_right_out[216]));

	mux_tree_tapbuf_size6 mux_right_track_440 (
		.in({chany_top_in[54], chany_top_in[128], chany_top_in[202], chany_top_in[276], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_36_sram_inv[0:2]),
		.out(chanx_right_out[220]));

	mux_tree_tapbuf_size6 mux_right_track_448 (
		.in({chany_top_in[55], chany_top_in[129], chany_top_in[203], chany_top_in[277], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_37_sram_inv[0:2]),
		.out(chanx_right_out[224]));

	mux_tree_tapbuf_size6 mux_right_track_456 (
		.in({chany_top_in[56], chany_top_in[130], chany_top_in[204], chany_top_in[278], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_38_sram_inv[0:2]),
		.out(chanx_right_out[228]));

	mux_tree_tapbuf_size6 mux_right_track_464 (
		.in({chany_top_in[57], chany_top_in[131], chany_top_in[205], chany_top_in[279], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_39_sram_inv[0:2]),
		.out(chanx_right_out[232]));

	mux_tree_tapbuf_size6 mux_right_track_472 (
		.in({chany_top_in[58], chany_top_in[132], chany_top_in[206], chany_top_in[280], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_40_sram_inv[0:2]),
		.out(chanx_right_out[236]));

	mux_tree_tapbuf_size6 mux_right_track_480 (
		.in({chany_top_in[59], chany_top_in[133], chany_top_in[207], chany_top_in[281], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_41_sram_inv[0:2]),
		.out(chanx_right_out[240]));

	mux_tree_tapbuf_size6 mux_right_track_504 (
		.in({chany_top_in[62], chany_top_in[136], chany_top_in[210], chany_top_in[284], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_42_sram_inv[0:2]),
		.out(chanx_right_out[252]));

	mux_tree_tapbuf_size6 mux_right_track_512 (
		.in({chany_top_in[63], chany_top_in[137], chany_top_in[211], chany_top_in[285], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_43_sram_inv[0:2]),
		.out(chanx_right_out[256]));

	mux_tree_tapbuf_size6 mux_right_track_520 (
		.in({chany_top_in[64], chany_top_in[138], chany_top_in[212], chany_top_in[286], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_44_sram_inv[0:2]),
		.out(chanx_right_out[260]));

	mux_tree_tapbuf_size6 mux_right_track_528 (
		.in({chany_top_in[65], chany_top_in[139], chany_top_in[213], chany_top_in[287], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_45_sram_inv[0:2]),
		.out(chanx_right_out[264]));

	mux_tree_tapbuf_size6 mux_right_track_536 (
		.in({chany_top_in[66], chany_top_in[140], chany_top_in[214], chany_top_in[288], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_46_sram_inv[0:2]),
		.out(chanx_right_out[268]));

	mux_tree_tapbuf_size6 mux_right_track_544 (
		.in({chany_top_in[67], chany_top_in[141], chany_top_in[215], chany_top_in[289], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_47_sram_inv[0:2]),
		.out(chanx_right_out[272]));

	mux_tree_tapbuf_size6 mux_right_track_552 (
		.in({chany_top_in[68], chany_top_in[142], chany_top_in[216], chany_top_in[290], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_48_sram_inv[0:2]),
		.out(chanx_right_out[276]));

	mux_tree_tapbuf_size6 mux_right_track_576 (
		.in({chany_top_in[71], chany_top_in[145], chany_top_in[219], chany_top_in[293], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_49_sram_inv[0:2]),
		.out(chanx_right_out[288]));

	mux_tree_tapbuf_size6 mux_right_track_584 (
		.in({chany_top_in[72], chany_top_in[146], chany_top_in[220], chany_top_in[294], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_50_sram_inv[0:2]),
		.out(chanx_right_out[292]));

	mux_tree_tapbuf_size6 mux_left_track_41 (
		.in({chany_top_in[69], chany_top_in[143], chany_top_in[217], chany_top_in[291], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_51_sram_inv[0:2]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size6 mux_left_track_49 (
		.in({chany_top_in[68], chany_top_in[142], chany_top_in[216], chany_top_in[290], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_52_sram_inv[0:2]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size6 mux_left_track_57 (
		.in({chany_top_in[67], chany_top_in[141], chany_top_in[215], chany_top_in[289], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_53_sram_inv[0:2]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size6 mux_left_track_65 (
		.in({chany_top_in[66], chany_top_in[140], chany_top_in[214], chany_top_in[288], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_54_sram_inv[0:2]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size6 mux_left_track_113 (
		.in({chany_top_in[60], chany_top_in[134], chany_top_in[208], chany_top_in[282], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_55_sram_inv[0:2]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size6 mux_left_track_121 (
		.in({chany_top_in[59], chany_top_in[133], chany_top_in[207], chany_top_in[281], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_56_sram_inv[0:2]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size6 mux_left_track_145 (
		.in({chany_top_in[56], chany_top_in[130], chany_top_in[204], chany_top_in[278], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_57_sram_inv[0:2]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size6 mux_left_track_153 (
		.in({chany_top_in[55], chany_top_in[129], chany_top_in[203], chany_top_in[277], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_58_sram_inv[0:2]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size6 mux_left_track_161 (
		.in({chany_top_in[54], chany_top_in[128], chany_top_in[202], chany_top_in[276], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_59_sram_inv[0:2]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size6 mux_left_track_169 (
		.in({chany_top_in[53], chany_top_in[127], chany_top_in[201], chany_top_in[275], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_60_sram_inv[0:2]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size6 mux_left_track_177 (
		.in({chany_top_in[52], chany_top_in[126], chany_top_in[200], chany_top_in[274], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_61_sram_inv[0:2]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size6 mux_left_track_185 (
		.in({chany_top_in[51], chany_top_in[125], chany_top_in[199], chany_top_in[273], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_62_sram_inv[0:2]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size6 mux_left_track_193 (
		.in({chany_top_in[50], chany_top_in[124], chany_top_in[198], chany_top_in[272], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_63_sram_inv[0:2]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size6 mux_left_track_217 (
		.in({chany_top_in[47], chany_top_in[121], chany_top_in[195], chany_top_in[269], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_64_sram_inv[0:2]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size6 mux_left_track_225 (
		.in({chany_top_in[46], chany_top_in[120], chany_top_in[194], chany_top_in[268], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_65_sram_inv[0:2]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size6 mux_left_track_233 (
		.in({chany_top_in[45], chany_top_in[119], chany_top_in[193], chany_top_in[267], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_66_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_66_sram_inv[0:2]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size6 mux_left_track_241 (
		.in({chany_top_in[44], chany_top_in[118], chany_top_in[192], chany_top_in[266], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_67_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_67_sram_inv[0:2]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size6 mux_left_track_249 (
		.in({chany_top_in[43], chany_top_in[117], chany_top_in[191], chany_top_in[265], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_68_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_68_sram_inv[0:2]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size6 mux_left_track_257 (
		.in({chany_top_in[42], chany_top_in[116], chany_top_in[190], chany_top_in[264], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_69_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_69_sram_inv[0:2]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size6 mux_left_track_265 (
		.in({chany_top_in[41], chany_top_in[115], chany_top_in[189], chany_top_in[263], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_70_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_70_sram_inv[0:2]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size6 mux_left_track_289 (
		.in({chany_top_in[38], chany_top_in[112], chany_top_in[186], chany_top_in[260], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_71_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_71_sram_inv[0:2]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size6 mux_left_track_297 (
		.in({chany_top_in[37], chany_top_in[111], chany_top_in[185], chany_top_in[259], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_72_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_72_sram_inv[0:2]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size6 mux_left_track_305 (
		.in({chany_top_in[36], chany_top_in[110], chany_top_in[184], chany_top_in[258], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_73_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_73_sram_inv[0:2]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size6 mux_left_track_313 (
		.in({chany_top_in[35], chany_top_in[109], chany_top_in[183], chany_top_in[257], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_74_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_74_sram_inv[0:2]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size6 mux_left_track_321 (
		.in({chany_top_in[34], chany_top_in[108], chany_top_in[182], chany_top_in[256], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_75_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_75_sram_inv[0:2]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size6 mux_left_track_329 (
		.in({chany_top_in[33], chany_top_in[107], chany_top_in[181], chany_top_in[255], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_76_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_76_sram_inv[0:2]),
		.out(chanx_left_out[164]));

	mux_tree_tapbuf_size6 mux_left_track_337 (
		.in({chany_top_in[32], chany_top_in[106], chany_top_in[180], chany_top_in[254], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_77_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_77_sram_inv[0:2]),
		.out(chanx_left_out[168]));

	mux_tree_tapbuf_size6 mux_left_track_361 (
		.in({chany_top_in[29], chany_top_in[103], chany_top_in[177], chany_top_in[251], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_78_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_78_sram_inv[0:2]),
		.out(chanx_left_out[180]));

	mux_tree_tapbuf_size6 mux_left_track_369 (
		.in({chany_top_in[28], chany_top_in[102], chany_top_in[176], chany_top_in[250], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_79_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_79_sram_inv[0:2]),
		.out(chanx_left_out[184]));

	mux_tree_tapbuf_size6 mux_left_track_377 (
		.in({chany_top_in[27], chany_top_in[101], chany_top_in[175], chany_top_in[249], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_80_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_80_sram_inv[0:2]),
		.out(chanx_left_out[188]));

	mux_tree_tapbuf_size6 mux_left_track_385 (
		.in({chany_top_in[26], chany_top_in[100], chany_top_in[174], chany_top_in[248], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_81_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_81_sram_inv[0:2]),
		.out(chanx_left_out[192]));

	mux_tree_tapbuf_size6 mux_left_track_393 (
		.in({chany_top_in[25], chany_top_in[99], chany_top_in[173], chany_top_in[247], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_82_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_82_sram_inv[0:2]),
		.out(chanx_left_out[196]));

	mux_tree_tapbuf_size6 mux_left_track_401 (
		.in({chany_top_in[24], chany_top_in[98], chany_top_in[172], chany_top_in[246], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_83_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_83_sram_inv[0:2]),
		.out(chanx_left_out[200]));

	mux_tree_tapbuf_size6 mux_left_track_409 (
		.in({chany_top_in[23], chany_top_in[97], chany_top_in[171], chany_top_in[245], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_84_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_84_sram_inv[0:2]),
		.out(chanx_left_out[204]));

	mux_tree_tapbuf_size6 mux_left_track_433 (
		.in({chany_top_in[20], chany_top_in[94], chany_top_in[168], chany_top_in[242], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_85_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_85_sram_inv[0:2]),
		.out(chanx_left_out[216]));

	mux_tree_tapbuf_size6 mux_left_track_441 (
		.in({chany_top_in[19], chany_top_in[93], chany_top_in[167], chany_top_in[241], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_86_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_86_sram_inv[0:2]),
		.out(chanx_left_out[220]));

	mux_tree_tapbuf_size6 mux_left_track_449 (
		.in({chany_top_in[18], chany_top_in[92], chany_top_in[166], chany_top_in[240], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_87_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_87_sram_inv[0:2]),
		.out(chanx_left_out[224]));

	mux_tree_tapbuf_size6 mux_left_track_457 (
		.in({chany_top_in[17], chany_top_in[91], chany_top_in[165], chany_top_in[239], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_88_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_88_sram_inv[0:2]),
		.out(chanx_left_out[228]));

	mux_tree_tapbuf_size6 mux_left_track_465 (
		.in({chany_top_in[16], chany_top_in[90], chany_top_in[164], chany_top_in[238], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_89_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_89_sram_inv[0:2]),
		.out(chanx_left_out[232]));

	mux_tree_tapbuf_size6 mux_left_track_473 (
		.in({chany_top_in[15], chany_top_in[89], chany_top_in[163], chany_top_in[237], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_90_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_90_sram_inv[0:2]),
		.out(chanx_left_out[236]));

	mux_tree_tapbuf_size6 mux_left_track_481 (
		.in({chany_top_in[14], chany_top_in[88], chany_top_in[162], chany_top_in[236], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_91_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_91_sram_inv[0:2]),
		.out(chanx_left_out[240]));

	mux_tree_tapbuf_size6 mux_left_track_505 (
		.in({chany_top_in[11], chany_top_in[85], chany_top_in[159], chany_top_in[233], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_92_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_92_sram_inv[0:2]),
		.out(chanx_left_out[252]));

	mux_tree_tapbuf_size6 mux_left_track_513 (
		.in({chany_top_in[10], chany_top_in[84], chany_top_in[158], chany_top_in[232], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_93_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_93_sram_inv[0:2]),
		.out(chanx_left_out[256]));

	mux_tree_tapbuf_size6 mux_left_track_521 (
		.in({chany_top_in[9], chany_top_in[83], chany_top_in[157], chany_top_in[231], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_94_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_94_sram_inv[0:2]),
		.out(chanx_left_out[260]));

	mux_tree_tapbuf_size6 mux_left_track_529 (
		.in({chany_top_in[8], chany_top_in[82], chany_top_in[156], chany_top_in[230], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_95_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_95_sram_inv[0:2]),
		.out(chanx_left_out[264]));

	mux_tree_tapbuf_size6 mux_left_track_537 (
		.in({chany_top_in[7], chany_top_in[81], chany_top_in[155], chany_top_in[229], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_96_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_96_sram_inv[0:2]),
		.out(chanx_left_out[268]));

	mux_tree_tapbuf_size6 mux_left_track_545 (
		.in({chany_top_in[6], chany_top_in[80], chany_top_in[154], chany_top_in[228], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_97_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_97_sram_inv[0:2]),
		.out(chanx_left_out[272]));

	mux_tree_tapbuf_size6 mux_left_track_553 (
		.in({chany_top_in[5], chany_top_in[79], chany_top_in[153], chany_top_in[227], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_98_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_98_sram_inv[0:2]),
		.out(chanx_left_out[276]));

	mux_tree_tapbuf_size6 mux_left_track_577 (
		.in({chany_top_in[2], chany_top_in[76], chany_top_in[150], chany_top_in[224], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_99_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_99_sram_inv[0:2]),
		.out(chanx_left_out[288]));

	mux_tree_tapbuf_size6 mux_left_track_585 (
		.in({chany_top_in[1], chany_top_in[75], chany_top_in[149], chany_top_in[223], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_100_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_100_sram_inv[0:2]),
		.out(chanx_left_out[292]));

	mux_tree_tapbuf_size6_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_11_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_12_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_13_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_14_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_15_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_16_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_17_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_18_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_19_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_20_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_21_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_22_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_23_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_24_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_25_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_26_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_27_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_28_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_29_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_30_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_31_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_32_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_33_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_34_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_35_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_36_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_37_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_38_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_39_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_40_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_41_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_42_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_43_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_44_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_45_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_46_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_47_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_48_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_576 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_49_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_584 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_50_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_51_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_52_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_53_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_54_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_55_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_56_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_57_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_58_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_59_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_60_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_61_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_62_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_63_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_64_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_65_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_66_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_66_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_67_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_67_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_68_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_68_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_69_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_69_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_70_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_70_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_71_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_71_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_72_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_72_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_73_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_73_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_74_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_74_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_75_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_75_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_76_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_76_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_77_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_77_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_78_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_78_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_79_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_79_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_80_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_80_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_81_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_81_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_393 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_82_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_82_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_401 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_83_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_83_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_409 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_84_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_84_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_433 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_85_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_85_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_441 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_86_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_86_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_449 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_87_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_87_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_457 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_88_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_88_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_465 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_89_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_89_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_473 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_90_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_90_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_481 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_91_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_91_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_505 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_92_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_92_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_513 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_93_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_93_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_521 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_94_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_94_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_529 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_95_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_95_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_537 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_96_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_96_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_545 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_97_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_97_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_553 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_98_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_98_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_577 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_99_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_99_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_585 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_99_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_100_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_100_sram_inv[0:2]));

	mux_tree_tapbuf_size4 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[2], chanx_right_in[11]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_size4 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[4], chanx_right_in[15]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_size4 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[5], chanx_right_in[19]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_size4 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[6], chanx_right_in[23]}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size4 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[8], chanx_right_in[27]}),
		.sram(mux_tree_tapbuf_size4_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_4_sram_inv[0:2]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_size4 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[9], chanx_right_in[31]}),
		.sram(mux_tree_tapbuf_size4_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_5_sram_inv[0:2]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_size4 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[10], chanx_right_in[35]}),
		.sram(mux_tree_tapbuf_size4_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_6_sram_inv[0:2]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_size4 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[13], chanx_right_in[43]}),
		.sram(mux_tree_tapbuf_size4_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_7_sram_inv[0:2]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_size4 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[14], chanx_right_in[47]}),
		.sram(mux_tree_tapbuf_size4_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_8_sram_inv[0:2]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_size4 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[16], chanx_right_in[51]}),
		.sram(mux_tree_tapbuf_size4_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_9_sram_inv[0:2]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_size4 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[17], chanx_right_in[55]}),
		.sram(mux_tree_tapbuf_size4_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_10_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size4 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[18], chanx_right_in[59]}),
		.sram(mux_tree_tapbuf_size4_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_11_sram_inv[0:2]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_size4 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[20], chanx_right_in[63]}),
		.sram(mux_tree_tapbuf_size4_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_12_sram_inv[0:2]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_size4 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[21], chanx_right_in[67]}),
		.sram(mux_tree_tapbuf_size4_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_13_sram_inv[0:2]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_size4 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[25], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size4_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_14_sram_inv[0:2]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_size4 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[26], chanx_right_in[83]}),
		.sram(mux_tree_tapbuf_size4_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_15_sram_inv[0:2]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_size4 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[28], chanx_right_in[87]}),
		.sram(mux_tree_tapbuf_size4_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_16_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size4 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[29], chanx_right_in[91]}),
		.sram(mux_tree_tapbuf_size4_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_17_sram_inv[0:2]),
		.out(chany_top_out[21]));

	mux_tree_tapbuf_size4 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[30], chanx_right_in[95]}),
		.sram(mux_tree_tapbuf_size4_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_18_sram_inv[0:2]),
		.out(chany_top_out[22]));

	mux_tree_tapbuf_size4 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[32], chanx_right_in[99]}),
		.sram(mux_tree_tapbuf_size4_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_19_sram_inv[0:2]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_size4 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[33], chanx_right_in[103]}),
		.sram(mux_tree_tapbuf_size4_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_20_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size4 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[37], chanx_right_in[115]}),
		.sram(mux_tree_tapbuf_size4_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_21_sram_inv[0:2]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_size4 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[38], chanx_right_in[119]}),
		.sram(mux_tree_tapbuf_size4_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_22_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size4 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[40], chanx_right_in[123]}),
		.sram(mux_tree_tapbuf_size4_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_23_sram_inv[0:2]),
		.out(chany_top_out[29]));

	mux_tree_tapbuf_size4 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[41], chanx_right_in[127]}),
		.sram(mux_tree_tapbuf_size4_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_24_sram_inv[0:2]),
		.out(chany_top_out[30]));

	mux_tree_tapbuf_size4 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[42], chanx_right_in[131]}),
		.sram(mux_tree_tapbuf_size4_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_25_sram_inv[0:2]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_size4 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[44], chanx_right_in[135]}),
		.sram(mux_tree_tapbuf_size4_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_26_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size4 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[45], chanx_right_in[139]}),
		.sram(mux_tree_tapbuf_size4_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_27_sram_inv[0:2]),
		.out(chany_top_out[33]));

	mux_tree_tapbuf_size4 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[49], chanx_right_in[151]}),
		.sram(mux_tree_tapbuf_size4_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_28_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size4 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[50], chanx_right_in[155]}),
		.sram(mux_tree_tapbuf_size4_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_29_sram_inv[0:2]),
		.out(chany_top_out[37]));

	mux_tree_tapbuf_size4 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[52], chanx_right_in[159]}),
		.sram(mux_tree_tapbuf_size4_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_30_sram_inv[0:2]),
		.out(chany_top_out[38]));

	mux_tree_tapbuf_size4 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[53], chanx_right_in[163]}),
		.sram(mux_tree_tapbuf_size4_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_31_sram_inv[0:2]),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_size4 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[54], chanx_right_in[167]}),
		.sram(mux_tree_tapbuf_size4_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_32_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size4 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[56], chanx_right_in[171]}),
		.sram(mux_tree_tapbuf_size4_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_33_sram_inv[0:2]),
		.out(chany_top_out[41]));

	mux_tree_tapbuf_size4 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[57], chanx_right_in[175]}),
		.sram(mux_tree_tapbuf_size4_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_34_sram_inv[0:2]),
		.out(chany_top_out[42]));

	mux_tree_tapbuf_size4 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[61], chanx_right_in[187]}),
		.sram(mux_tree_tapbuf_size4_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_35_sram_inv[0:2]),
		.out(chany_top_out[45]));

	mux_tree_tapbuf_size4 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[62], chanx_right_in[191]}),
		.sram(mux_tree_tapbuf_size4_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_36_sram_inv[0:2]),
		.out(chany_top_out[46]));

	mux_tree_tapbuf_size4 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[64], chanx_right_in[195]}),
		.sram(mux_tree_tapbuf_size4_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_37_sram_inv[0:2]),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_size4 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[65], chanx_right_in[199]}),
		.sram(mux_tree_tapbuf_size4_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_38_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size4 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[66], chanx_right_in[203]}),
		.sram(mux_tree_tapbuf_size4_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_39_sram_inv[0:2]),
		.out(chany_top_out[49]));

	mux_tree_tapbuf_size4 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[68], chanx_right_in[207]}),
		.sram(mux_tree_tapbuf_size4_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_40_sram_inv[0:2]),
		.out(chany_top_out[50]));

	mux_tree_tapbuf_size4 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[69], chanx_right_in[211]}),
		.sram(mux_tree_tapbuf_size4_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_41_sram_inv[0:2]),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_size4 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[73], chanx_right_in[223]}),
		.sram(mux_tree_tapbuf_size4_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_42_sram_inv[0:2]),
		.out(chany_top_out[54]));

	mux_tree_tapbuf_size4 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[74], chanx_right_in[227]}),
		.sram(mux_tree_tapbuf_size4_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_43_sram_inv[0:2]),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_size4 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[76], chanx_right_in[231]}),
		.sram(mux_tree_tapbuf_size4_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_44_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size4 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[77], chanx_right_in[235]}),
		.sram(mux_tree_tapbuf_size4_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_45_sram_inv[0:2]),
		.out(chany_top_out[57]));

	mux_tree_tapbuf_size4 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[78], chanx_right_in[239]}),
		.sram(mux_tree_tapbuf_size4_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_46_sram_inv[0:2]),
		.out(chany_top_out[58]));

	mux_tree_tapbuf_size4 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[80], chanx_right_in[243]}),
		.sram(mux_tree_tapbuf_size4_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_47_sram_inv[0:2]),
		.out(chany_top_out[59]));

	mux_tree_tapbuf_size4 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[81], chanx_right_in[247]}),
		.sram(mux_tree_tapbuf_size4_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_48_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size4 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[85], chanx_right_in[259]}),
		.sram(mux_tree_tapbuf_size4_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_49_sram_inv[0:2]),
		.out(chany_top_out[63]));

	mux_tree_tapbuf_size4 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[86], chanx_right_in[263]}),
		.sram(mux_tree_tapbuf_size4_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_50_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size4 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[88], chanx_right_in[267]}),
		.sram(mux_tree_tapbuf_size4_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_51_sram_inv[0:2]),
		.out(chany_top_out[65]));

	mux_tree_tapbuf_size4 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[89], chanx_right_in[271]}),
		.sram(mux_tree_tapbuf_size4_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_52_sram_inv[0:2]),
		.out(chany_top_out[66]));

	mux_tree_tapbuf_size4 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[90], chanx_right_in[275]}),
		.sram(mux_tree_tapbuf_size4_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_53_sram_inv[0:2]),
		.out(chany_top_out[67]));

	mux_tree_tapbuf_size4 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[92], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size4_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_54_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size4 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[93], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size4_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_55_sram_inv[0:2]),
		.out(chany_top_out[69]));

	mux_tree_tapbuf_size4 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[97], chanx_right_in[295]}),
		.sram(mux_tree_tapbuf_size4_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_56_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size4 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[101], chanx_left_in[294]}),
		.sram(mux_tree_tapbuf_size4_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_57_sram_inv[0:2]),
		.out(chany_top_out[75]));

	mux_tree_tapbuf_size4 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[102], chanx_left_in[293]}),
		.sram(mux_tree_tapbuf_size4_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_58_sram_inv[0:2]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size4 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[104], chanx_left_in[292]}),
		.sram(mux_tree_tapbuf_size4_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_59_sram_inv[0:2]),
		.out(chany_top_out[77]));

	mux_tree_tapbuf_size4 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[105], chanx_left_in[290]}),
		.sram(mux_tree_tapbuf_size4_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_60_sram_inv[0:2]),
		.out(chany_top_out[78]));

	mux_tree_tapbuf_size4 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[109], chanx_left_in[286]}),
		.sram(mux_tree_tapbuf_size4_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_61_sram_inv[0:2]),
		.out(chany_top_out[81]));

	mux_tree_tapbuf_size4 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[110], chanx_left_in[285]}),
		.sram(mux_tree_tapbuf_size4_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_62_sram_inv[0:2]),
		.out(chany_top_out[82]));

	mux_tree_tapbuf_size4 mux_top_track_166 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[112], chanx_left_in[284]}),
		.sram(mux_tree_tapbuf_size4_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_63_sram_inv[0:2]),
		.out(chany_top_out[83]));

	mux_tree_tapbuf_size4 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[113], chanx_left_in[282]}),
		.sram(mux_tree_tapbuf_size4_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_64_sram_inv[0:2]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size4 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[114], chanx_left_in[281]}),
		.sram(mux_tree_tapbuf_size4_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_65_sram_inv[0:2]),
		.out(chany_top_out[85]));

	mux_tree_tapbuf_size4 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[116], chanx_left_in[280]}),
		.sram(mux_tree_tapbuf_size4_66_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_66_sram_inv[0:2]),
		.out(chany_top_out[86]));

	mux_tree_tapbuf_size4 mux_top_track_174 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[117], chanx_left_in[278]}),
		.sram(mux_tree_tapbuf_size4_67_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_67_sram_inv[0:2]),
		.out(chany_top_out[87]));

	mux_tree_tapbuf_size4 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[121], chanx_left_in[274]}),
		.sram(mux_tree_tapbuf_size4_68_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_68_sram_inv[0:2]),
		.out(chany_top_out[90]));

	mux_tree_tapbuf_size4 mux_top_track_182 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[122], chanx_left_in[273]}),
		.sram(mux_tree_tapbuf_size4_69_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_69_sram_inv[0:2]),
		.out(chany_top_out[91]));

	mux_tree_tapbuf_size4 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[124], chanx_left_in[272]}),
		.sram(mux_tree_tapbuf_size4_70_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_70_sram_inv[0:2]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size4 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[125], chanx_left_in[270]}),
		.sram(mux_tree_tapbuf_size4_71_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_71_sram_inv[0:2]),
		.out(chany_top_out[93]));

	mux_tree_tapbuf_size4 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[126], chanx_left_in[269]}),
		.sram(mux_tree_tapbuf_size4_72_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_72_sram_inv[0:2]),
		.out(chany_top_out[94]));

	mux_tree_tapbuf_size4 mux_top_track_190 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[128], chanx_left_in[268]}),
		.sram(mux_tree_tapbuf_size4_73_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_73_sram_inv[0:2]),
		.out(chany_top_out[95]));

	mux_tree_tapbuf_size4 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[129], chanx_left_in[266]}),
		.sram(mux_tree_tapbuf_size4_74_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_74_sram_inv[0:2]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size4 mux_top_track_198 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[133], chanx_left_in[262]}),
		.sram(mux_tree_tapbuf_size4_75_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_75_sram_inv[0:2]),
		.out(chany_top_out[99]));

	mux_tree_tapbuf_size4 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[134], chanx_left_in[261]}),
		.sram(mux_tree_tapbuf_size4_76_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_76_sram_inv[0:2]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size4 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[136], chanx_left_in[260]}),
		.sram(mux_tree_tapbuf_size4_77_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_77_sram_inv[0:2]),
		.out(chany_top_out[101]));

	mux_tree_tapbuf_size4 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[137], chanx_left_in[258]}),
		.sram(mux_tree_tapbuf_size4_78_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_78_sram_inv[0:2]),
		.out(chany_top_out[102]));

	mux_tree_tapbuf_size4 mux_top_track_206 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[138], chanx_left_in[257]}),
		.sram(mux_tree_tapbuf_size4_79_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_79_sram_inv[0:2]),
		.out(chany_top_out[103]));

	mux_tree_tapbuf_size4 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[140], chanx_left_in[256]}),
		.sram(mux_tree_tapbuf_size4_80_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_80_sram_inv[0:2]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size4 mux_top_track_210 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[141], chanx_left_in[254]}),
		.sram(mux_tree_tapbuf_size4_81_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_81_sram_inv[0:2]),
		.out(chany_top_out[105]));

	mux_tree_tapbuf_size4 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[145], chanx_left_in[250]}),
		.sram(mux_tree_tapbuf_size4_82_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_82_sram_inv[0:2]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size4 mux_top_track_218 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[146], chanx_left_in[249]}),
		.sram(mux_tree_tapbuf_size4_83_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_83_sram_inv[0:2]),
		.out(chany_top_out[109]));

	mux_tree_tapbuf_size4 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[148], chanx_left_in[248]}),
		.sram(mux_tree_tapbuf_size4_84_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_84_sram_inv[0:2]),
		.out(chany_top_out[110]));

	mux_tree_tapbuf_size4 mux_top_track_222 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[149], chanx_left_in[246]}),
		.sram(mux_tree_tapbuf_size4_85_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_85_sram_inv[0:2]),
		.out(chany_top_out[111]));

	mux_tree_tapbuf_size4 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[150], chanx_left_in[245]}),
		.sram(mux_tree_tapbuf_size4_86_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_86_sram_inv[0:2]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size4 mux_top_track_226 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[152], chanx_left_in[244]}),
		.sram(mux_tree_tapbuf_size4_87_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_87_sram_inv[0:2]),
		.out(chany_top_out[113]));

	mux_tree_tapbuf_size4 mux_top_track_228 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[153], chanx_left_in[242]}),
		.sram(mux_tree_tapbuf_size4_88_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_88_sram_inv[0:2]),
		.out(chany_top_out[114]));

	mux_tree_tapbuf_size4 mux_top_track_234 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[157], chanx_left_in[238]}),
		.sram(mux_tree_tapbuf_size4_89_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_89_sram_inv[0:2]),
		.out(chany_top_out[117]));

	mux_tree_tapbuf_size4 mux_top_track_236 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[158], chanx_left_in[237]}),
		.sram(mux_tree_tapbuf_size4_90_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_90_sram_inv[0:2]),
		.out(chany_top_out[118]));

	mux_tree_tapbuf_size4 mux_top_track_238 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[160], chanx_left_in[236]}),
		.sram(mux_tree_tapbuf_size4_91_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_91_sram_inv[0:2]),
		.out(chany_top_out[119]));

	mux_tree_tapbuf_size4 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[161], chanx_left_in[234]}),
		.sram(mux_tree_tapbuf_size4_92_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_92_sram_inv[0:2]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size4 mux_top_track_242 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[162], chanx_left_in[233]}),
		.sram(mux_tree_tapbuf_size4_93_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_93_sram_inv[0:2]),
		.out(chany_top_out[121]));

	mux_tree_tapbuf_size4 mux_top_track_244 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[164], chanx_left_in[232]}),
		.sram(mux_tree_tapbuf_size4_94_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_94_sram_inv[0:2]),
		.out(chany_top_out[122]));

	mux_tree_tapbuf_size4 mux_top_track_246 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[165], chanx_left_in[230]}),
		.sram(mux_tree_tapbuf_size4_95_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_95_sram_inv[0:2]),
		.out(chany_top_out[123]));

	mux_tree_tapbuf_size4 mux_top_track_252 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[169], chanx_left_in[226]}),
		.sram(mux_tree_tapbuf_size4_96_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_96_sram_inv[0:2]),
		.out(chany_top_out[126]));

	mux_tree_tapbuf_size4 mux_top_track_254 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[170], chanx_left_in[225]}),
		.sram(mux_tree_tapbuf_size4_97_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_97_sram_inv[0:2]),
		.out(chany_top_out[127]));

	mux_tree_tapbuf_size4 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[172], chanx_left_in[224]}),
		.sram(mux_tree_tapbuf_size4_98_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_98_sram_inv[0:2]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size4 mux_top_track_258 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[173], chanx_left_in[222]}),
		.sram(mux_tree_tapbuf_size4_99_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_99_sram_inv[0:2]),
		.out(chany_top_out[129]));

	mux_tree_tapbuf_size4 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[174], chanx_left_in[221]}),
		.sram(mux_tree_tapbuf_size4_100_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_100_sram_inv[0:2]),
		.out(chany_top_out[130]));

	mux_tree_tapbuf_size4 mux_top_track_262 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[176], chanx_left_in[220]}),
		.sram(mux_tree_tapbuf_size4_101_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_101_sram_inv[0:2]),
		.out(chany_top_out[131]));

	mux_tree_tapbuf_size4 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[177], chanx_left_in[218]}),
		.sram(mux_tree_tapbuf_size4_102_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_102_sram_inv[0:2]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size4 mux_top_track_270 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[181], chanx_left_in[214]}),
		.sram(mux_tree_tapbuf_size4_103_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_103_sram_inv[0:2]),
		.out(chany_top_out[135]));

	mux_tree_tapbuf_size4 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[182], chanx_left_in[213]}),
		.sram(mux_tree_tapbuf_size4_104_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_104_sram_inv[0:2]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size4 mux_top_track_274 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[184], chanx_left_in[212]}),
		.sram(mux_tree_tapbuf_size4_105_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_105_sram_inv[0:2]),
		.out(chany_top_out[137]));

	mux_tree_tapbuf_size4 mux_top_track_276 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[185], chanx_left_in[210]}),
		.sram(mux_tree_tapbuf_size4_106_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_106_sram_inv[0:2]),
		.out(chany_top_out[138]));

	mux_tree_tapbuf_size4 mux_top_track_278 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[186], chanx_left_in[209]}),
		.sram(mux_tree_tapbuf_size4_107_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_107_sram_inv[0:2]),
		.out(chany_top_out[139]));

	mux_tree_tapbuf_size4 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[188], chanx_left_in[208]}),
		.sram(mux_tree_tapbuf_size4_108_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_108_sram_inv[0:2]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size4 mux_top_track_282 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[189], chanx_left_in[206]}),
		.sram(mux_tree_tapbuf_size4_109_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_109_sram_inv[0:2]),
		.out(chany_top_out[141]));

	mux_tree_tapbuf_size4 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[193], chanx_left_in[202]}),
		.sram(mux_tree_tapbuf_size4_110_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_110_sram_inv[0:2]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size4 mux_top_track_290 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[194], chanx_left_in[201]}),
		.sram(mux_tree_tapbuf_size4_111_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_111_sram_inv[0:2]),
		.out(chany_top_out[145]));

	mux_tree_tapbuf_size4 mux_top_track_292 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[196], chanx_left_in[200]}),
		.sram(mux_tree_tapbuf_size4_112_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_112_sram_inv[0:2]),
		.out(chany_top_out[146]));

	mux_tree_tapbuf_size4 mux_top_track_294 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[197], chanx_left_in[198]}),
		.sram(mux_tree_tapbuf_size4_113_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_113_sram_inv[0:2]),
		.out(chany_top_out[147]));

	mux_tree_tapbuf_size4 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[198], chanx_left_in[197]}),
		.sram(mux_tree_tapbuf_size4_114_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_114_sram_inv[0:2]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size4 mux_top_track_298 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[200], chanx_left_in[196]}),
		.sram(mux_tree_tapbuf_size4_115_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_115_sram_inv[0:2]),
		.out(chany_top_out[149]));

	mux_tree_tapbuf_size4 mux_top_track_300 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[201], chanx_left_in[194]}),
		.sram(mux_tree_tapbuf_size4_116_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_116_sram_inv[0:2]),
		.out(chany_top_out[150]));

	mux_tree_tapbuf_size4 mux_top_track_306 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[205], chanx_left_in[190]}),
		.sram(mux_tree_tapbuf_size4_117_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_117_sram_inv[0:2]),
		.out(chany_top_out[153]));

	mux_tree_tapbuf_size4 mux_top_track_308 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[206], chanx_left_in[189]}),
		.sram(mux_tree_tapbuf_size4_118_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_118_sram_inv[0:2]),
		.out(chany_top_out[154]));

	mux_tree_tapbuf_size4 mux_top_track_310 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[208], chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size4_119_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_119_sram_inv[0:2]),
		.out(chany_top_out[155]));

	mux_tree_tapbuf_size4 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[209], chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size4_120_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_120_sram_inv[0:2]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size4 mux_top_track_314 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[210], chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size4_121_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_121_sram_inv[0:2]),
		.out(chany_top_out[157]));

	mux_tree_tapbuf_size4 mux_top_track_316 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[212], chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size4_122_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_122_sram_inv[0:2]),
		.out(chany_top_out[158]));

	mux_tree_tapbuf_size4 mux_top_track_318 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[213], chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size4_123_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_123_sram_inv[0:2]),
		.out(chany_top_out[159]));

	mux_tree_tapbuf_size4 mux_top_track_324 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[217], chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size4_124_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_124_sram_inv[0:2]),
		.out(chany_top_out[162]));

	mux_tree_tapbuf_size4 mux_top_track_326 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[218], chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size4_125_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_125_sram_inv[0:2]),
		.out(chany_top_out[163]));

	mux_tree_tapbuf_size4 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[220], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size4_126_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_126_sram_inv[0:2]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size4 mux_top_track_330 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[221], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size4_127_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_127_sram_inv[0:2]),
		.out(chany_top_out[165]));

	mux_tree_tapbuf_size4 mux_top_track_332 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[222], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size4_128_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_128_sram_inv[0:2]),
		.out(chany_top_out[166]));

	mux_tree_tapbuf_size4 mux_top_track_334 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[224], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size4_129_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_129_sram_inv[0:2]),
		.out(chany_top_out[167]));

	mux_tree_tapbuf_size4 mux_top_track_336 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[225], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size4_130_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_130_sram_inv[0:2]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size4 mux_top_track_342 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[229], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size4_131_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_131_sram_inv[0:2]),
		.out(chany_top_out[171]));

	mux_tree_tapbuf_size4 mux_top_track_344 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[230], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size4_132_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_132_sram_inv[0:2]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size4 mux_top_track_346 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[232], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size4_133_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_133_sram_inv[0:2]),
		.out(chany_top_out[173]));

	mux_tree_tapbuf_size4 mux_top_track_348 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[233], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size4_134_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_134_sram_inv[0:2]),
		.out(chany_top_out[174]));

	mux_tree_tapbuf_size4 mux_top_track_350 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[234], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size4_135_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_135_sram_inv[0:2]),
		.out(chany_top_out[175]));

	mux_tree_tapbuf_size4 mux_top_track_352 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[236], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size4_136_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_136_sram_inv[0:2]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size4 mux_top_track_354 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[237], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size4_137_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_137_sram_inv[0:2]),
		.out(chany_top_out[177]));

	mux_tree_tapbuf_size4 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[241], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size4_138_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_138_sram_inv[0:2]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size4 mux_top_track_362 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[242], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size4_139_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_139_sram_inv[0:2]),
		.out(chany_top_out[181]));

	mux_tree_tapbuf_size4 mux_top_track_364 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[244], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size4_140_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_140_sram_inv[0:2]),
		.out(chany_top_out[182]));

	mux_tree_tapbuf_size4 mux_top_track_366 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[245], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size4_141_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_141_sram_inv[0:2]),
		.out(chany_top_out[183]));

	mux_tree_tapbuf_size4 mux_top_track_368 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[246], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size4_142_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_142_sram_inv[0:2]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size4 mux_top_track_370 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[248], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size4_143_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_143_sram_inv[0:2]),
		.out(chany_top_out[185]));

	mux_tree_tapbuf_size4 mux_top_track_372 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[249], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size4_144_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_144_sram_inv[0:2]),
		.out(chany_top_out[186]));

	mux_tree_tapbuf_size4 mux_top_track_378 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[253], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size4_145_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_145_sram_inv[0:2]),
		.out(chany_top_out[189]));

	mux_tree_tapbuf_size4 mux_top_track_380 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[254], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size4_146_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_146_sram_inv[0:2]),
		.out(chany_top_out[190]));

	mux_tree_tapbuf_size4 mux_top_track_382 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[256], chanx_left_in[140]}),
		.sram(mux_tree_tapbuf_size4_147_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_147_sram_inv[0:2]),
		.out(chany_top_out[191]));

	mux_tree_tapbuf_size4 mux_top_track_384 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[257], chanx_left_in[138]}),
		.sram(mux_tree_tapbuf_size4_148_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_148_sram_inv[0:2]),
		.out(chany_top_out[192]));

	mux_tree_tapbuf_size4 mux_top_track_386 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[258], chanx_left_in[137]}),
		.sram(mux_tree_tapbuf_size4_149_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_149_sram_inv[0:2]),
		.out(chany_top_out[193]));

	mux_tree_tapbuf_size4 mux_top_track_388 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[260], chanx_left_in[136]}),
		.sram(mux_tree_tapbuf_size4_150_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_150_sram_inv[0:2]),
		.out(chany_top_out[194]));

	mux_tree_tapbuf_size4 mux_top_track_390 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[261], chanx_left_in[134]}),
		.sram(mux_tree_tapbuf_size4_151_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_151_sram_inv[0:2]),
		.out(chany_top_out[195]));

	mux_tree_tapbuf_size4 mux_top_track_396 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[265], chanx_left_in[130]}),
		.sram(mux_tree_tapbuf_size4_152_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_152_sram_inv[0:2]),
		.out(chany_top_out[198]));

	mux_tree_tapbuf_size4 mux_top_track_398 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[266], chanx_left_in[129]}),
		.sram(mux_tree_tapbuf_size4_153_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_153_sram_inv[0:2]),
		.out(chany_top_out[199]));

	mux_tree_tapbuf_size4 mux_top_track_400 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[268], chanx_left_in[128]}),
		.sram(mux_tree_tapbuf_size4_154_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_154_sram_inv[0:2]),
		.out(chany_top_out[200]));

	mux_tree_tapbuf_size4 mux_top_track_402 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[269], chanx_left_in[126]}),
		.sram(mux_tree_tapbuf_size4_155_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_155_sram_inv[0:2]),
		.out(chany_top_out[201]));

	mux_tree_tapbuf_size4 mux_top_track_404 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[270], chanx_left_in[125]}),
		.sram(mux_tree_tapbuf_size4_156_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_156_sram_inv[0:2]),
		.out(chany_top_out[202]));

	mux_tree_tapbuf_size4 mux_top_track_406 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[272], chanx_left_in[124]}),
		.sram(mux_tree_tapbuf_size4_157_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_157_sram_inv[0:2]),
		.out(chany_top_out[203]));

	mux_tree_tapbuf_size4 mux_top_track_408 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[273], chanx_left_in[122]}),
		.sram(mux_tree_tapbuf_size4_158_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_158_sram_inv[0:2]),
		.out(chany_top_out[204]));

	mux_tree_tapbuf_size4 mux_top_track_414 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[277], chanx_left_in[118]}),
		.sram(mux_tree_tapbuf_size4_159_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_159_sram_inv[0:2]),
		.out(chany_top_out[207]));

	mux_tree_tapbuf_size4 mux_top_track_416 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[278], chanx_left_in[117]}),
		.sram(mux_tree_tapbuf_size4_160_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_160_sram_inv[0:2]),
		.out(chany_top_out[208]));

	mux_tree_tapbuf_size4 mux_top_track_418 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[280], chanx_left_in[116]}),
		.sram(mux_tree_tapbuf_size4_161_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_161_sram_inv[0:2]),
		.out(chany_top_out[209]));

	mux_tree_tapbuf_size4 mux_top_track_420 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[281], chanx_left_in[114]}),
		.sram(mux_tree_tapbuf_size4_162_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_162_sram_inv[0:2]),
		.out(chany_top_out[210]));

	mux_tree_tapbuf_size4 mux_top_track_422 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[282], chanx_left_in[113]}),
		.sram(mux_tree_tapbuf_size4_163_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_163_sram_inv[0:2]),
		.out(chany_top_out[211]));

	mux_tree_tapbuf_size4 mux_top_track_424 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[284], chanx_left_in[112]}),
		.sram(mux_tree_tapbuf_size4_164_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_164_sram_inv[0:2]),
		.out(chany_top_out[212]));

	mux_tree_tapbuf_size4 mux_top_track_426 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[285], chanx_left_in[110]}),
		.sram(mux_tree_tapbuf_size4_165_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_165_sram_inv[0:2]),
		.out(chany_top_out[213]));

	mux_tree_tapbuf_size4 mux_top_track_432 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[289], chanx_left_in[106]}),
		.sram(mux_tree_tapbuf_size4_166_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_166_sram_inv[0:2]),
		.out(chany_top_out[216]));

	mux_tree_tapbuf_size4 mux_top_track_434 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[290], chanx_left_in[105]}),
		.sram(mux_tree_tapbuf_size4_167_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_167_sram_inv[0:2]),
		.out(chany_top_out[217]));

	mux_tree_tapbuf_size4 mux_top_track_436 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[292], chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size4_168_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_168_sram_inv[0:2]),
		.out(chany_top_out[218]));

	mux_tree_tapbuf_size4 mux_top_track_438 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[293], chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size4_169_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_169_sram_inv[0:2]),
		.out(chany_top_out[219]));

	mux_tree_tapbuf_size4 mux_top_track_440 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[294], chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size4_170_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_170_sram_inv[0:2]),
		.out(chany_top_out[220]));

	mux_tree_tapbuf_size4 mux_top_track_450 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[94], chanx_left_in[287]}),
		.sram(mux_tree_tapbuf_size4_171_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_171_sram_inv[0:2]),
		.out(chany_top_out[225]));

	mux_tree_tapbuf_size4 mux_top_track_452 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[93], chanx_left_in[283]}),
		.sram(mux_tree_tapbuf_size4_172_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_172_sram_inv[0:2]),
		.out(chany_top_out[226]));

	mux_tree_tapbuf_size4 mux_top_track_454 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[92], chanx_left_in[279]}),
		.sram(mux_tree_tapbuf_size4_173_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_173_sram_inv[0:2]),
		.out(chany_top_out[227]));

	mux_tree_tapbuf_size4 mux_top_track_456 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[90], chanx_left_in[275]}),
		.sram(mux_tree_tapbuf_size4_174_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_174_sram_inv[0:2]),
		.out(chany_top_out[228]));

	mux_tree_tapbuf_size4 mux_top_track_458 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[89], chanx_left_in[271]}),
		.sram(mux_tree_tapbuf_size4_175_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_175_sram_inv[0:2]),
		.out(chany_top_out[229]));

	mux_tree_tapbuf_size4 mux_top_track_460 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[88], chanx_left_in[267]}),
		.sram(mux_tree_tapbuf_size4_176_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_176_sram_inv[0:2]),
		.out(chany_top_out[230]));

	mux_tree_tapbuf_size4 mux_top_track_462 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[86], chanx_left_in[263]}),
		.sram(mux_tree_tapbuf_size4_177_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_177_sram_inv[0:2]),
		.out(chany_top_out[231]));

	mux_tree_tapbuf_size4 mux_top_track_468 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[82], chanx_left_in[251]}),
		.sram(mux_tree_tapbuf_size4_178_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_178_sram_inv[0:2]),
		.out(chany_top_out[234]));

	mux_tree_tapbuf_size4 mux_top_track_470 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[81], chanx_left_in[247]}),
		.sram(mux_tree_tapbuf_size4_179_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_179_sram_inv[0:2]),
		.out(chany_top_out[235]));

	mux_tree_tapbuf_size4 mux_top_track_472 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[80], chanx_left_in[243]}),
		.sram(mux_tree_tapbuf_size4_180_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_180_sram_inv[0:2]),
		.out(chany_top_out[236]));

	mux_tree_tapbuf_size4 mux_top_track_474 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[78], chanx_left_in[239]}),
		.sram(mux_tree_tapbuf_size4_181_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_181_sram_inv[0:2]),
		.out(chany_top_out[237]));

	mux_tree_tapbuf_size4 mux_top_track_476 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[77], chanx_left_in[235]}),
		.sram(mux_tree_tapbuf_size4_182_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_182_sram_inv[0:2]),
		.out(chany_top_out[238]));

	mux_tree_tapbuf_size4 mux_top_track_478 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[76], chanx_left_in[231]}),
		.sram(mux_tree_tapbuf_size4_183_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_183_sram_inv[0:2]),
		.out(chany_top_out[239]));

	mux_tree_tapbuf_size4 mux_top_track_480 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[74], chanx_left_in[227]}),
		.sram(mux_tree_tapbuf_size4_184_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_184_sram_inv[0:2]),
		.out(chany_top_out[240]));

	mux_tree_tapbuf_size4 mux_top_track_486 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[70], chanx_left_in[215]}),
		.sram(mux_tree_tapbuf_size4_185_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_185_sram_inv[0:2]),
		.out(chany_top_out[243]));

	mux_tree_tapbuf_size4 mux_top_track_488 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[69], chanx_left_in[211]}),
		.sram(mux_tree_tapbuf_size4_186_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_186_sram_inv[0:2]),
		.out(chany_top_out[244]));

	mux_tree_tapbuf_size4 mux_top_track_490 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[68], chanx_left_in[207]}),
		.sram(mux_tree_tapbuf_size4_187_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_187_sram_inv[0:2]),
		.out(chany_top_out[245]));

	mux_tree_tapbuf_size4 mux_top_track_492 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[66], chanx_left_in[203]}),
		.sram(mux_tree_tapbuf_size4_188_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_188_sram_inv[0:2]),
		.out(chany_top_out[246]));

	mux_tree_tapbuf_size4 mux_top_track_494 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[65], chanx_left_in[199]}),
		.sram(mux_tree_tapbuf_size4_189_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_189_sram_inv[0:2]),
		.out(chany_top_out[247]));

	mux_tree_tapbuf_size4 mux_top_track_496 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[64], chanx_left_in[195]}),
		.sram(mux_tree_tapbuf_size4_190_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_190_sram_inv[0:2]),
		.out(chany_top_out[248]));

	mux_tree_tapbuf_size4 mux_top_track_498 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[62], chanx_left_in[191]}),
		.sram(mux_tree_tapbuf_size4_191_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_191_sram_inv[0:2]),
		.out(chany_top_out[249]));

	mux_tree_tapbuf_size4 mux_top_track_504 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[58], chanx_left_in[179]}),
		.sram(mux_tree_tapbuf_size4_192_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_192_sram_inv[0:2]),
		.out(chany_top_out[252]));

	mux_tree_tapbuf_size4 mux_top_track_506 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[57], chanx_left_in[175]}),
		.sram(mux_tree_tapbuf_size4_193_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_193_sram_inv[0:2]),
		.out(chany_top_out[253]));

	mux_tree_tapbuf_size4 mux_top_track_508 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[56], chanx_left_in[171]}),
		.sram(mux_tree_tapbuf_size4_194_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_194_sram_inv[0:2]),
		.out(chany_top_out[254]));

	mux_tree_tapbuf_size4 mux_top_track_510 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[54], chanx_left_in[167]}),
		.sram(mux_tree_tapbuf_size4_195_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_195_sram_inv[0:2]),
		.out(chany_top_out[255]));

	mux_tree_tapbuf_size4 mux_top_track_512 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[53], chanx_left_in[163]}),
		.sram(mux_tree_tapbuf_size4_196_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_196_sram_inv[0:2]),
		.out(chany_top_out[256]));

	mux_tree_tapbuf_size4 mux_top_track_514 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[52], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size4_197_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_197_sram_inv[0:2]),
		.out(chany_top_out[257]));

	mux_tree_tapbuf_size4 mux_top_track_516 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[50], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size4_198_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_198_sram_inv[0:2]),
		.out(chany_top_out[258]));

	mux_tree_tapbuf_size4 mux_top_track_522 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[46], chanx_left_in[143]}),
		.sram(mux_tree_tapbuf_size4_199_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_199_sram_inv[0:2]),
		.out(chany_top_out[261]));

	mux_tree_tapbuf_size4 mux_top_track_524 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[45], chanx_left_in[139]}),
		.sram(mux_tree_tapbuf_size4_200_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_200_sram_inv[0:2]),
		.out(chany_top_out[262]));

	mux_tree_tapbuf_size4 mux_top_track_526 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[44], chanx_left_in[135]}),
		.sram(mux_tree_tapbuf_size4_201_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_201_sram_inv[0:2]),
		.out(chany_top_out[263]));

	mux_tree_tapbuf_size4 mux_top_track_528 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[42], chanx_left_in[131]}),
		.sram(mux_tree_tapbuf_size4_202_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_202_sram_inv[0:2]),
		.out(chany_top_out[264]));

	mux_tree_tapbuf_size4 mux_top_track_530 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[41], chanx_left_in[127]}),
		.sram(mux_tree_tapbuf_size4_203_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_203_sram_inv[0:2]),
		.out(chany_top_out[265]));

	mux_tree_tapbuf_size4 mux_top_track_532 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[40], chanx_left_in[123]}),
		.sram(mux_tree_tapbuf_size4_204_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_204_sram_inv[0:2]),
		.out(chany_top_out[266]));

	mux_tree_tapbuf_size4 mux_top_track_534 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[38], chanx_left_in[119]}),
		.sram(mux_tree_tapbuf_size4_205_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_205_sram_inv[0:2]),
		.out(chany_top_out[267]));

	mux_tree_tapbuf_size4 mux_top_track_540 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[34], chanx_left_in[107]}),
		.sram(mux_tree_tapbuf_size4_206_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_206_sram_inv[0:2]),
		.out(chany_top_out[270]));

	mux_tree_tapbuf_size4 mux_top_track_542 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[33], chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size4_207_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_207_sram_inv[0:2]),
		.out(chany_top_out[271]));

	mux_tree_tapbuf_size4 mux_top_track_544 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[32], chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size4_208_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_208_sram_inv[0:2]),
		.out(chany_top_out[272]));

	mux_tree_tapbuf_size4 mux_top_track_546 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[30], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_size4_209_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_209_sram_inv[0:2]),
		.out(chany_top_out[273]));

	mux_tree_tapbuf_size4 mux_top_track_548 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[29], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_size4_210_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_210_sram_inv[0:2]),
		.out(chany_top_out[274]));

	mux_tree_tapbuf_size4 mux_top_track_550 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[28], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_size4_211_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_211_sram_inv[0:2]),
		.out(chany_top_out[275]));

	mux_tree_tapbuf_size4 mux_top_track_552 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[26], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_size4_212_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_212_sram_inv[0:2]),
		.out(chany_top_out[276]));

	mux_tree_tapbuf_size4 mux_top_track_558 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[22], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_size4_213_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_213_sram_inv[0:2]),
		.out(chany_top_out[279]));

	mux_tree_tapbuf_size4 mux_top_track_560 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[21], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_size4_214_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_214_sram_inv[0:2]),
		.out(chany_top_out[280]));

	mux_tree_tapbuf_size4 mux_top_track_562 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[20], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_size4_215_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_215_sram_inv[0:2]),
		.out(chany_top_out[281]));

	mux_tree_tapbuf_size4 mux_top_track_564 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[18], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_size4_216_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_216_sram_inv[0:2]),
		.out(chany_top_out[282]));

	mux_tree_tapbuf_size4 mux_top_track_566 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[17], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_size4_217_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_217_sram_inv[0:2]),
		.out(chany_top_out[283]));

	mux_tree_tapbuf_size4 mux_top_track_568 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[16], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_size4_218_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_218_sram_inv[0:2]),
		.out(chany_top_out[284]));

	mux_tree_tapbuf_size4 mux_top_track_570 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[14], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_size4_219_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_219_sram_inv[0:2]),
		.out(chany_top_out[285]));

	mux_tree_tapbuf_size4 mux_top_track_576 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[10], chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_size4_220_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_220_sram_inv[0:2]),
		.out(chany_top_out[288]));

	mux_tree_tapbuf_size4 mux_top_track_578 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[9], chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_size4_221_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_221_sram_inv[0:2]),
		.out(chany_top_out[289]));

	mux_tree_tapbuf_size4 mux_top_track_580 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[8], chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_size4_222_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_222_sram_inv[0:2]),
		.out(chany_top_out[290]));

	mux_tree_tapbuf_size4 mux_top_track_582 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[6], chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_size4_223_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_223_sram_inv[0:2]),
		.out(chany_top_out[291]));

	mux_tree_tapbuf_size4 mux_top_track_584 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[5], chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_size4_224_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_224_sram_inv[0:2]),
		.out(chany_top_out[292]));

	mux_tree_tapbuf_size4 mux_top_track_586 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[4], chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_size4_225_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_225_sram_inv[0:2]),
		.out(chany_top_out[293]));

	mux_tree_tapbuf_size4 mux_top_track_588 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[2], chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_size4_226_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_226_sram_inv[0:2]),
		.out(chany_top_out[294]));

	mux_tree_tapbuf_size4_mem mem_top_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_4_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_5_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_6_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_7_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_8_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_9_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_10_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_11_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_12_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_13_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_14_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_15_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_16_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_17_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_18_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_19_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_20_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_21_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_22_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_23_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_24_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_25_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_26_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_27_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_28_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_29_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_30_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_31_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_32_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_33_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_34_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_35_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_36_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_37_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_38_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_39_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_40_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_41_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_42_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_43_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_44_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_45_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_46_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_47_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_48_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_49_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_50_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_51_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_52_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_53_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_54_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_55_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_56_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_57_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_58_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_59_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_60_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_61_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_62_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_63_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_64_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_65_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_66_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_66_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_67_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_67_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_68_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_68_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_69_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_69_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_70_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_70_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_71_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_71_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_72_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_72_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_73_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_73_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_74_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_74_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_75_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_75_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_76_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_76_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_77_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_77_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_78_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_78_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_79_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_79_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_80_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_80_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_81_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_81_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_82_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_82_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_218 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_83_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_83_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_220 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_84_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_84_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_222 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_85_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_85_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_86_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_86_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_226 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_87_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_87_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_228 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_88_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_88_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_234 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_89_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_89_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_236 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_90_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_90_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_238 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_91_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_91_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_92_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_92_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_242 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_93_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_93_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_244 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_94_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_94_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_246 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_95_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_95_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_252 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_96_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_96_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_254 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_97_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_97_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_98_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_98_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_258 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_99_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_99_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_260 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_100_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_100_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_262 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_101_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_101_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_102_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_102_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_270 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_103_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_103_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_104_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_104_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_274 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_105_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_105_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_276 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_106_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_106_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_278 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_107_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_107_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_108_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_108_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_282 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_109_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_109_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_110_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_110_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_290 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_111_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_111_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_292 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_112_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_112_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_294 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_113_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_113_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_114_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_114_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_298 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_115_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_115_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_300 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_116_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_116_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_306 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_117_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_117_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_308 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_118_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_118_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_310 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_119_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_119_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_120_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_120_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_314 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_121_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_121_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_316 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_122_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_122_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_318 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_123_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_123_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_324 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_124_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_124_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_326 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_125_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_125_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_126_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_126_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_330 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_127_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_127_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_332 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_128_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_128_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_334 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_129_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_129_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_130_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_130_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_342 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_131_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_131_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_132_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_132_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_346 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_133_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_133_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_348 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_134_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_134_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_350 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_135_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_135_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_136_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_136_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_136_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_354 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_136_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_137_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_137_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_137_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_138_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_138_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_138_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_362 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_138_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_139_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_139_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_139_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_364 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_139_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_140_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_140_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_140_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_366 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_140_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_141_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_141_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_141_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_141_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_142_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_142_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_142_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_370 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_142_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_143_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_143_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_143_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_372 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_143_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_144_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_144_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_144_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_378 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_145_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_145_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_145_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_380 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_145_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_146_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_146_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_146_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_382 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_146_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_147_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_147_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_147_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_147_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_148_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_148_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_148_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_386 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_148_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_149_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_149_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_149_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_388 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_149_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_150_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_150_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_150_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_390 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_150_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_151_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_151_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_151_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_396 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_152_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_152_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_152_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_398 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_152_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_153_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_153_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_153_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_153_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_154_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_154_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_154_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_402 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_154_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_155_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_155_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_155_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_404 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_155_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_156_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_156_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_156_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_406 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_156_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_157_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_157_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_157_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_157_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_158_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_158_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_158_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_414 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_159_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_159_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_159_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_159_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_160_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_160_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_160_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_418 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_160_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_161_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_161_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_161_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_420 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_161_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_162_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_162_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_162_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_422 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_162_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_163_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_163_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_163_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_163_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_164_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_164_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_164_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_426 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_164_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_165_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_165_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_165_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_166_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_166_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_166_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_434 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_166_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_167_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_167_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_167_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_436 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_167_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_168_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_168_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_168_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_438 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_168_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_169_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_169_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_169_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_169_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_170_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_170_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_170_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_450 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_171_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_171_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_171_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_452 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_171_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_172_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_172_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_172_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_454 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_172_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_173_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_173_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_173_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_173_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_174_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_174_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_174_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_458 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_174_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_175_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_175_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_175_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_460 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_175_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_176_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_176_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_176_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_462 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_176_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_177_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_177_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_177_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_468 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_178_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_178_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_178_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_470 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_178_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_179_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_179_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_179_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_179_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_180_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_180_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_180_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_474 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_180_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_181_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_181_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_181_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_476 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_181_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_182_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_182_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_182_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_478 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_182_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_183_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_183_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_183_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_183_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_184_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_184_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_184_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_486 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_185_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_185_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_185_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_185_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_186_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_186_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_186_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_490 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_186_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_187_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_187_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_187_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_492 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_187_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_188_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_188_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_188_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_494 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_188_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_189_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_189_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_189_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_189_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_190_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_190_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_190_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_498 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_190_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_191_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_191_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_191_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_192_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_192_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_192_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_506 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_192_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_193_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_193_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_193_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_508 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_193_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_194_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_194_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_194_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_510 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_194_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_195_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_195_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_195_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_195_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_196_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_196_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_196_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_514 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_196_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_197_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_197_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_197_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_516 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_197_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_198_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_198_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_198_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_522 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_199_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_199_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_199_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_524 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_199_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_200_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_200_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_200_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_526 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_200_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_201_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_201_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_201_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_201_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_202_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_202_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_202_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_530 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_202_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_203_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_203_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_203_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_532 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_203_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_204_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_204_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_204_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_534 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_204_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_205_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_205_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_205_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_540 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_206_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_206_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_206_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_542 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_206_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_207_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_207_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_207_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_207_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_208_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_208_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_208_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_546 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_208_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_209_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_209_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_209_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_548 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_209_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_210_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_210_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_210_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_550 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_210_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_211_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_211_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_211_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_211_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_212_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_212_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_212_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_558 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_213_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_213_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_213_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_213_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_214_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_214_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_214_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_562 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_214_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_215_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_215_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_215_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_564 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_215_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_216_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_216_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_216_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_566 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_216_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_217_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_217_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_217_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_217_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_218_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_218_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_218_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_570 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_218_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_219_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_219_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_219_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_576 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_220_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_220_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_220_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_578 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_220_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_221_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_221_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_221_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_580 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_221_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_222_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_222_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_222_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_582 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_222_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_223_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_223_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_223_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_584 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_223_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_224_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_224_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_224_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_586 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_224_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_225_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_225_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_225_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_588 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_225_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_226_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_226_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_226_sram_inv[0:2]));

	mux_tree_tapbuf_size3 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[12], chanx_right_in[39]}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size3 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[22], chanx_right_in[71]}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size3 mux_top_track_34 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[24], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_size3 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[34], chanx_right_in[107]}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_tree_tapbuf_size3 mux_top_track_52 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[36], chanx_right_in[111]}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chany_top_out[26]));

	mux_tree_tapbuf_size3 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[46], chanx_right_in[143]}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_tree_tapbuf_size3 mux_top_track_70 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[48], chanx_right_in[147]}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_size3 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[58], chanx_right_in[179]}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_size3 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[60], chanx_right_in[183]}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size3 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[70], chanx_right_in[215]}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size3 mux_top_track_106 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[72], chanx_right_in[219]}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chany_top_out[53]));

	mux_tree_tapbuf_size3 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[82], chanx_right_in[251]}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chany_top_out[61]));

	mux_tree_tapbuf_size3 mux_top_track_124 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[84], chanx_right_in[255]}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chany_top_out[62]));

	mux_tree_tapbuf_size3 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[94], chanx_right_in[287]}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chany_top_out[70]));

	mux_tree_tapbuf_size3 mux_top_track_142 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[96], chanx_right_in[291]}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chany_top_out[71]));

	mux_tree_tapbuf_size3 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[98]}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_tree_tapbuf_size3 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[100]}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_tree_tapbuf_size3 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[106], chanx_left_in[289]}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_tree_tapbuf_size3 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[108], chanx_left_in[288]}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size3 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[118], chanx_left_in[277]}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size3 mux_top_track_178 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[120], chanx_left_in[276]}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_top_out[89]));

	mux_tree_tapbuf_size3 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[130], chanx_left_in[265]}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_top_out[97]));

	mux_tree_tapbuf_size3 mux_top_track_196 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[132], chanx_left_in[264]}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_top_out[98]));

	mux_tree_tapbuf_size3 mux_top_track_212 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[142], chanx_left_in[253]}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_top_out[106]));

	mux_tree_tapbuf_size3 mux_top_track_214 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[144], chanx_left_in[252]}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_top_out[107]));

	mux_tree_tapbuf_size3 mux_top_track_230 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[154], chanx_left_in[241]}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_top_out[115]));

	mux_tree_tapbuf_size3 mux_top_track_232 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[156], chanx_left_in[240]}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size3 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[166], chanx_left_in[229]}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size3 mux_top_track_250 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[168], chanx_left_in[228]}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_top_out[125]));

	mux_tree_tapbuf_size3 mux_top_track_266 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[178], chanx_left_in[217]}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_top_out[133]));

	mux_tree_tapbuf_size3 mux_top_track_268 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[180], chanx_left_in[216]}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chany_top_out[134]));

	mux_tree_tapbuf_size3 mux_top_track_284 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[190], chanx_left_in[205]}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chany_top_out[142]));

	mux_tree_tapbuf_size3 mux_top_track_286 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[192], chanx_left_in[204]}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chany_top_out[143]));

	mux_tree_tapbuf_size3 mux_top_track_302 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[202], chanx_left_in[193]}),
		.sram(mux_tree_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_33_sram_inv[0:1]),
		.out(chany_top_out[151]));

	mux_tree_tapbuf_size3 mux_top_track_304 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[204], chanx_left_in[192]}),
		.sram(mux_tree_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_34_sram_inv[0:1]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size3 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[214], chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_35_sram_inv[0:1]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size3 mux_top_track_322 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[216], chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_36_sram_inv[0:1]),
		.out(chany_top_out[161]));

	mux_tree_tapbuf_size3 mux_top_track_338 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[226], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_37_sram_inv[0:1]),
		.out(chany_top_out[169]));

	mux_tree_tapbuf_size3 mux_top_track_340 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[228], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_38_sram_inv[0:1]),
		.out(chany_top_out[170]));

	mux_tree_tapbuf_size3 mux_top_track_356 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[238], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_39_sram_inv[0:1]),
		.out(chany_top_out[178]));

	mux_tree_tapbuf_size3 mux_top_track_358 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[240], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_40_sram_inv[0:1]),
		.out(chany_top_out[179]));

	mux_tree_tapbuf_size3 mux_top_track_374 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[250], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_41_sram_inv[0:1]),
		.out(chany_top_out[187]));

	mux_tree_tapbuf_size3 mux_top_track_376 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[252], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_42_sram_inv[0:1]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size3 mux_top_track_392 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[262], chanx_left_in[133]}),
		.sram(mux_tree_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_43_sram_inv[0:1]),
		.out(chany_top_out[196]));

	mux_tree_tapbuf_size3 mux_top_track_394 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[264], chanx_left_in[132]}),
		.sram(mux_tree_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_44_sram_inv[0:1]),
		.out(chany_top_out[197]));

	mux_tree_tapbuf_size3 mux_top_track_410 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[274], chanx_left_in[121]}),
		.sram(mux_tree_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_45_sram_inv[0:1]),
		.out(chany_top_out[205]));

	mux_tree_tapbuf_size3 mux_top_track_412 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[276], chanx_left_in[120]}),
		.sram(mux_tree_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_46_sram_inv[0:1]),
		.out(chany_top_out[206]));

	mux_tree_tapbuf_size3 mux_top_track_428 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[286], chanx_left_in[109]}),
		.sram(mux_tree_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_47_sram_inv[0:1]),
		.out(chany_top_out[214]));

	mux_tree_tapbuf_size3 mux_top_track_430 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[288], chanx_left_in[108]}),
		.sram(mux_tree_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_48_sram_inv[0:1]),
		.out(chany_top_out[215]));

	mux_tree_tapbuf_size3 mux_top_track_442 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_49_sram_inv[0:1]),
		.out(chany_top_out[221]));

	mux_tree_tapbuf_size3 mux_top_track_444 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_50_sram_inv[0:1]),
		.out(chany_top_out[222]));

	mux_tree_tapbuf_size3 mux_top_track_446 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[97], chanx_left_in[295]}),
		.sram(mux_tree_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_51_sram_inv[0:1]),
		.out(chany_top_out[223]));

	mux_tree_tapbuf_size3 mux_top_track_448 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[96], chanx_left_in[291]}),
		.sram(mux_tree_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_52_sram_inv[0:1]),
		.out(chany_top_out[224]));

	mux_tree_tapbuf_size3 mux_top_track_464 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[85], chanx_left_in[259]}),
		.sram(mux_tree_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_53_sram_inv[0:1]),
		.out(chany_top_out[232]));

	mux_tree_tapbuf_size3 mux_top_track_466 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[84], chanx_left_in[255]}),
		.sram(mux_tree_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_54_sram_inv[0:1]),
		.out(chany_top_out[233]));

	mux_tree_tapbuf_size3 mux_top_track_482 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[73], chanx_left_in[223]}),
		.sram(mux_tree_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_55_sram_inv[0:1]),
		.out(chany_top_out[241]));

	mux_tree_tapbuf_size3 mux_top_track_484 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[72], chanx_left_in[219]}),
		.sram(mux_tree_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_56_sram_inv[0:1]),
		.out(chany_top_out[242]));

	mux_tree_tapbuf_size3 mux_top_track_500 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[61], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_57_sram_inv[0:1]),
		.out(chany_top_out[250]));

	mux_tree_tapbuf_size3 mux_top_track_502 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[60], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_58_sram_inv[0:1]),
		.out(chany_top_out[251]));

	mux_tree_tapbuf_size3 mux_top_track_518 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[49], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_59_sram_inv[0:1]),
		.out(chany_top_out[259]));

	mux_tree_tapbuf_size3 mux_top_track_520 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[48], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_60_sram_inv[0:1]),
		.out(chany_top_out[260]));

	mux_tree_tapbuf_size3 mux_top_track_536 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[37], chanx_left_in[115]}),
		.sram(mux_tree_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_61_sram_inv[0:1]),
		.out(chany_top_out[268]));

	mux_tree_tapbuf_size3 mux_top_track_538 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[36], chanx_left_in[111]}),
		.sram(mux_tree_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_62_sram_inv[0:1]),
		.out(chany_top_out[269]));

	mux_tree_tapbuf_size3 mux_top_track_554 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[25], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_63_sram_inv[0:1]),
		.out(chany_top_out[277]));

	mux_tree_tapbuf_size3 mux_top_track_556 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[24], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_64_sram_inv[0:1]),
		.out(chany_top_out[278]));

	mux_tree_tapbuf_size3 mux_top_track_572 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[13], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_65_sram_inv[0:1]),
		.out(chany_top_out[286]));

	mux_tree_tapbuf_size3 mux_top_track_574 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[12], chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_66_sram_inv[0:1]),
		.out(chany_top_out[287]));

	mux_tree_tapbuf_size3_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_212 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_214 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_230 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_250 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_266 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_268 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_284 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_286 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_302 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_322 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_338 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_340 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_356 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_137_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_358 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_374 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_144_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_151_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_394 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_410 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_158_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_412 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_428 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_165_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_430 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_442 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_170_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_444 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_446 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_177_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_466 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_482 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_184_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_55_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_484 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_56_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_500 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_191_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_57_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_502 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_58_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_518 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_198_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_59_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_60_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_205_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_61_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_538 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_62_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_554 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_212_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_63_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_556 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_64_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_572 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_219_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_65_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_574 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_66_sram_inv[0:1]));

	mux_tree_tapbuf_size5 mux_top_track_590 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[0], chanx_right_in[3], chanx_left_in[1], chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_top_out[295]));

	mux_tree_tapbuf_size5 mux_right_track_128 (
		.in({chany_top_in[15], chany_top_in[89], chany_top_in[163], chany_top_in[237], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size5 mux_right_track_136 (
		.in({chany_top_in[16], chany_top_in[90], chany_top_in[164], chany_top_in[238], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size5 mux_right_track_200 (
		.in({chany_top_in[24], chany_top_in[98], chany_top_in[172], chany_top_in[246], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size5 mux_right_track_208 (
		.in({chany_top_in[25], chany_top_in[99], chany_top_in[173], chany_top_in[247], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size5 mux_right_track_272 (
		.in({chany_top_in[33], chany_top_in[107], chany_top_in[181], chany_top_in[255], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size5 mux_right_track_280 (
		.in({chany_top_in[34], chany_top_in[108], chany_top_in[182], chany_top_in[256], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size5 mux_right_track_344 (
		.in({chany_top_in[42], chany_top_in[116], chany_top_in[190], chany_top_in[264], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size5 mux_right_track_352 (
		.in({chany_top_in[43], chany_top_in[117], chany_top_in[191], chany_top_in[265], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size5 mux_right_track_416 (
		.in({chany_top_in[51], chany_top_in[125], chany_top_in[199], chany_top_in[273], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chanx_right_out[208]));

	mux_tree_tapbuf_size5 mux_right_track_424 (
		.in({chany_top_in[52], chany_top_in[126], chany_top_in[200], chany_top_in[274], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chanx_right_out[212]));

	mux_tree_tapbuf_size5 mux_right_track_488 (
		.in({chany_top_in[60], chany_top_in[134], chany_top_in[208], chany_top_in[282], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chanx_right_out[244]));

	mux_tree_tapbuf_size5 mux_right_track_496 (
		.in({chany_top_in[61], chany_top_in[135], chany_top_in[209], chany_top_in[283], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chanx_right_out[248]));

	mux_tree_tapbuf_size5 mux_right_track_560 (
		.in({chany_top_in[69], chany_top_in[143], chany_top_in[217], chany_top_in[291], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chanx_right_out[280]));

	mux_tree_tapbuf_size5 mux_right_track_568 (
		.in({chany_top_in[70], chany_top_in[144], chany_top_in[218], chany_top_in[292], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chanx_right_out[284]));

	mux_tree_tapbuf_size5 mux_left_track_129 (
		.in({chany_top_in[58], chany_top_in[132], chany_top_in[206], chany_top_in[280], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size5 mux_left_track_137 (
		.in({chany_top_in[57], chany_top_in[131], chany_top_in[205], chany_top_in[279], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size5 mux_left_track_201 (
		.in({chany_top_in[49], chany_top_in[123], chany_top_in[197], chany_top_in[271], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size5 mux_left_track_209 (
		.in({chany_top_in[48], chany_top_in[122], chany_top_in[196], chany_top_in[270], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size5 mux_left_track_273 (
		.in({chany_top_in[40], chany_top_in[114], chany_top_in[188], chany_top_in[262], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size5 mux_left_track_281 (
		.in({chany_top_in[39], chany_top_in[113], chany_top_in[187], chany_top_in[261], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size5 mux_left_track_345 (
		.in({chany_top_in[31], chany_top_in[105], chany_top_in[179], chany_top_in[253], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chanx_left_out[172]));

	mux_tree_tapbuf_size5 mux_left_track_353 (
		.in({chany_top_in[30], chany_top_in[104], chany_top_in[178], chany_top_in[252], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chanx_left_out[176]));

	mux_tree_tapbuf_size5 mux_left_track_417 (
		.in({chany_top_in[22], chany_top_in[96], chany_top_in[170], chany_top_in[244], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chanx_left_out[208]));

	mux_tree_tapbuf_size5 mux_left_track_425 (
		.in({chany_top_in[21], chany_top_in[95], chany_top_in[169], chany_top_in[243], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chanx_left_out[212]));

	mux_tree_tapbuf_size5 mux_left_track_489 (
		.in({chany_top_in[13], chany_top_in[87], chany_top_in[161], chany_top_in[235], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chanx_left_out[244]));

	mux_tree_tapbuf_size5 mux_left_track_497 (
		.in({chany_top_in[12], chany_top_in[86], chany_top_in[160], chany_top_in[234], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chanx_left_out[248]));

	mux_tree_tapbuf_size5 mux_left_track_561 (
		.in({chany_top_in[4], chany_top_in[78], chany_top_in[152], chany_top_in[226], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chanx_left_out[280]));

	mux_tree_tapbuf_size5 mux_left_track_569 (
		.in({chany_top_in[3], chany_top_in[77], chany_top_in[151], chany_top_in[225], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chanx_left_out[284]));

	mux_tree_tapbuf_size5_mem mem_top_track_590 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_226_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_417 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_425 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_489 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_497 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_561 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_569 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size7 mux_right_track_0 (
		.in({chany_top_in[73], chany_top_in[147], chany_top_in[221], chany_top_in[295], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size7 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[74], chany_top_in[148], chany_top_in[222], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size7 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[75], chany_top_in[149], chany_top_in[223], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size7 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[76], chany_top_in[150], chany_top_in[224], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_3_sram_inv[0:2]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size7 mux_right_track_32 (
		.in({chany_top_in[3], chany_top_in[77], chany_top_in[151], chany_top_in[225], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_4_sram_inv[0:2]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size7 mux_right_track_72 (
		.in({chany_top_in[8], chany_top_in[82], chany_top_in[156], chany_top_in[230], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_5_sram_inv[0:2]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size7 mux_right_track_80 (
		.in({chany_top_in[9], chany_top_in[83], chany_top_in[157], chany_top_in[231], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_6_sram_inv[0:2]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size7 mux_right_track_88 (
		.in({chany_top_in[10], chany_top_in[84], chany_top_in[158], chany_top_in[232], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_7_sram_inv[0:2]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size7 mux_right_track_96 (
		.in({chany_top_in[11], chany_top_in[85], chany_top_in[159], chany_top_in[233], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_8_sram_inv[0:2]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size7 mux_right_track_104 (
		.in({chany_top_in[12], chany_top_in[86], chany_top_in[160], chany_top_in[234], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_9_sram_inv[0:2]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size7 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[74], chany_top_in[148], chany_top_in[222], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_10_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size7 mux_left_track_9 (
		.in({chany_top_in[73], chany_top_in[147], chany_top_in[221], chany_top_in[295], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_11_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size7 mux_left_track_17 (
		.in({chany_top_in[72], chany_top_in[146], chany_top_in[220], chany_top_in[294], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_12_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size7 mux_left_track_25 (
		.in({chany_top_in[71], chany_top_in[145], chany_top_in[219], chany_top_in[293], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_13_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size7 mux_left_track_33 (
		.in({chany_top_in[70], chany_top_in[144], chany_top_in[218], chany_top_in[292], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_14_sram_inv[0:2]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size7 mux_left_track_73 (
		.in({chany_top_in[65], chany_top_in[139], chany_top_in[213], chany_top_in[287], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_15_sram_inv[0:2]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size7 mux_left_track_81 (
		.in({chany_top_in[64], chany_top_in[138], chany_top_in[212], chany_top_in[286], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_16_sram_inv[0:2]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size7 mux_left_track_89 (
		.in({chany_top_in[63], chany_top_in[137], chany_top_in[211], chany_top_in[285], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_17_sram_inv[0:2]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size7 mux_left_track_97 (
		.in({chany_top_in[62], chany_top_in[136], chany_top_in[210], chany_top_in[284], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_18_sram_inv[0:2]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size7 mux_left_track_105 (
		.in({chany_top_in[61], chany_top_in[135], chany_top_in[209], chany_top_in[283], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_19_sram_inv[0:2]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size7_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_9_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_10_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_11_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_12_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_13_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_14_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_15_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_16_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_17_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_18_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_19_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_1__0_ -----

//----- Default net type -----
`default_nettype wire



