//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jun 28 13:25:01 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_1__0_ -----
module sb_1__0_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:176] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:176] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:176] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:176] chany_top_out;
//----- OUTPUT PORTS -----
output [0:176] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:176] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_100_sram;
wire [0:1] mux_tree_tapbuf_size2_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_101_sram;
wire [0:1] mux_tree_tapbuf_size2_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_102_sram;
wire [0:1] mux_tree_tapbuf_size2_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_103_sram;
wire [0:1] mux_tree_tapbuf_size2_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_104_sram;
wire [0:1] mux_tree_tapbuf_size2_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_105_sram;
wire [0:1] mux_tree_tapbuf_size2_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_106_sram;
wire [0:1] mux_tree_tapbuf_size2_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_107_sram;
wire [0:1] mux_tree_tapbuf_size2_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_108_sram;
wire [0:1] mux_tree_tapbuf_size2_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_109_sram;
wire [0:1] mux_tree_tapbuf_size2_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_110_sram;
wire [0:1] mux_tree_tapbuf_size2_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_111_sram;
wire [0:1] mux_tree_tapbuf_size2_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_112_sram;
wire [0:1] mux_tree_tapbuf_size2_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_113_sram;
wire [0:1] mux_tree_tapbuf_size2_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_114_sram;
wire [0:1] mux_tree_tapbuf_size2_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_115_sram;
wire [0:1] mux_tree_tapbuf_size2_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_116_sram;
wire [0:1] mux_tree_tapbuf_size2_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_117_sram;
wire [0:1] mux_tree_tapbuf_size2_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_118_sram;
wire [0:1] mux_tree_tapbuf_size2_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_119_sram;
wire [0:1] mux_tree_tapbuf_size2_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_120_sram;
wire [0:1] mux_tree_tapbuf_size2_120_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_121_sram;
wire [0:1] mux_tree_tapbuf_size2_121_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_122_sram;
wire [0:1] mux_tree_tapbuf_size2_122_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_123_sram;
wire [0:1] mux_tree_tapbuf_size2_123_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_124_sram;
wire [0:1] mux_tree_tapbuf_size2_124_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_125_sram;
wire [0:1] mux_tree_tapbuf_size2_125_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_126_sram;
wire [0:1] mux_tree_tapbuf_size2_126_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_127_sram;
wire [0:1] mux_tree_tapbuf_size2_127_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_128_sram;
wire [0:1] mux_tree_tapbuf_size2_128_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_129_sram;
wire [0:1] mux_tree_tapbuf_size2_129_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_130_sram;
wire [0:1] mux_tree_tapbuf_size2_130_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_131_sram;
wire [0:1] mux_tree_tapbuf_size2_131_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_132_sram;
wire [0:1] mux_tree_tapbuf_size2_132_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_133_sram;
wire [0:1] mux_tree_tapbuf_size2_133_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_134_sram;
wire [0:1] mux_tree_tapbuf_size2_134_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_135_sram;
wire [0:1] mux_tree_tapbuf_size2_135_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_16_sram;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_17_sram;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_18_sram;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_19_sram;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_20_sram;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_21_sram;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_22_sram;
wire [0:1] mux_tree_tapbuf_size2_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_23_sram;
wire [0:1] mux_tree_tapbuf_size2_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_24_sram;
wire [0:1] mux_tree_tapbuf_size2_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_25_sram;
wire [0:1] mux_tree_tapbuf_size2_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_26_sram;
wire [0:1] mux_tree_tapbuf_size2_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_27_sram;
wire [0:1] mux_tree_tapbuf_size2_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_28_sram;
wire [0:1] mux_tree_tapbuf_size2_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_29_sram;
wire [0:1] mux_tree_tapbuf_size2_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_30_sram;
wire [0:1] mux_tree_tapbuf_size2_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_31_sram;
wire [0:1] mux_tree_tapbuf_size2_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_32_sram;
wire [0:1] mux_tree_tapbuf_size2_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_33_sram;
wire [0:1] mux_tree_tapbuf_size2_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_34_sram;
wire [0:1] mux_tree_tapbuf_size2_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_35_sram;
wire [0:1] mux_tree_tapbuf_size2_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_36_sram;
wire [0:1] mux_tree_tapbuf_size2_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_37_sram;
wire [0:1] mux_tree_tapbuf_size2_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_38_sram;
wire [0:1] mux_tree_tapbuf_size2_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_39_sram;
wire [0:1] mux_tree_tapbuf_size2_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_40_sram;
wire [0:1] mux_tree_tapbuf_size2_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_41_sram;
wire [0:1] mux_tree_tapbuf_size2_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_42_sram;
wire [0:1] mux_tree_tapbuf_size2_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_43_sram;
wire [0:1] mux_tree_tapbuf_size2_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_44_sram;
wire [0:1] mux_tree_tapbuf_size2_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_45_sram;
wire [0:1] mux_tree_tapbuf_size2_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_46_sram;
wire [0:1] mux_tree_tapbuf_size2_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_47_sram;
wire [0:1] mux_tree_tapbuf_size2_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_48_sram;
wire [0:1] mux_tree_tapbuf_size2_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_49_sram;
wire [0:1] mux_tree_tapbuf_size2_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_50_sram;
wire [0:1] mux_tree_tapbuf_size2_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_51_sram;
wire [0:1] mux_tree_tapbuf_size2_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_52_sram;
wire [0:1] mux_tree_tapbuf_size2_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_53_sram;
wire [0:1] mux_tree_tapbuf_size2_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_54_sram;
wire [0:1] mux_tree_tapbuf_size2_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_55_sram;
wire [0:1] mux_tree_tapbuf_size2_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_56_sram;
wire [0:1] mux_tree_tapbuf_size2_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_57_sram;
wire [0:1] mux_tree_tapbuf_size2_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_58_sram;
wire [0:1] mux_tree_tapbuf_size2_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_59_sram;
wire [0:1] mux_tree_tapbuf_size2_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_60_sram;
wire [0:1] mux_tree_tapbuf_size2_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_61_sram;
wire [0:1] mux_tree_tapbuf_size2_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_62_sram;
wire [0:1] mux_tree_tapbuf_size2_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_63_sram;
wire [0:1] mux_tree_tapbuf_size2_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_64_sram;
wire [0:1] mux_tree_tapbuf_size2_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_65_sram;
wire [0:1] mux_tree_tapbuf_size2_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_66_sram;
wire [0:1] mux_tree_tapbuf_size2_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_67_sram;
wire [0:1] mux_tree_tapbuf_size2_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_68_sram;
wire [0:1] mux_tree_tapbuf_size2_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_69_sram;
wire [0:1] mux_tree_tapbuf_size2_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_70_sram;
wire [0:1] mux_tree_tapbuf_size2_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_71_sram;
wire [0:1] mux_tree_tapbuf_size2_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_72_sram;
wire [0:1] mux_tree_tapbuf_size2_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_73_sram;
wire [0:1] mux_tree_tapbuf_size2_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_74_sram;
wire [0:1] mux_tree_tapbuf_size2_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_75_sram;
wire [0:1] mux_tree_tapbuf_size2_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_76_sram;
wire [0:1] mux_tree_tapbuf_size2_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_77_sram;
wire [0:1] mux_tree_tapbuf_size2_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_78_sram;
wire [0:1] mux_tree_tapbuf_size2_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_79_sram;
wire [0:1] mux_tree_tapbuf_size2_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_80_sram;
wire [0:1] mux_tree_tapbuf_size2_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_81_sram;
wire [0:1] mux_tree_tapbuf_size2_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_82_sram;
wire [0:1] mux_tree_tapbuf_size2_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_83_sram;
wire [0:1] mux_tree_tapbuf_size2_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_84_sram;
wire [0:1] mux_tree_tapbuf_size2_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_85_sram;
wire [0:1] mux_tree_tapbuf_size2_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_86_sram;
wire [0:1] mux_tree_tapbuf_size2_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_87_sram;
wire [0:1] mux_tree_tapbuf_size2_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_88_sram;
wire [0:1] mux_tree_tapbuf_size2_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_89_sram;
wire [0:1] mux_tree_tapbuf_size2_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_90_sram;
wire [0:1] mux_tree_tapbuf_size2_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_91_sram;
wire [0:1] mux_tree_tapbuf_size2_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_92_sram;
wire [0:1] mux_tree_tapbuf_size2_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_93_sram;
wire [0:1] mux_tree_tapbuf_size2_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_94_sram;
wire [0:1] mux_tree_tapbuf_size2_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_95_sram;
wire [0:1] mux_tree_tapbuf_size2_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_96_sram;
wire [0:1] mux_tree_tapbuf_size2_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_97_sram;
wire [0:1] mux_tree_tapbuf_size2_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_98_sram;
wire [0:1] mux_tree_tapbuf_size2_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_99_sram;
wire [0:1] mux_tree_tapbuf_size2_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_4_sram;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_5_sram;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_6_sram;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_7_sram;
wire [0:2] mux_tree_tapbuf_size4_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_8_sram;
wire [0:2] mux_tree_tapbuf_size4_8_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_8_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_29_sram;
wire [0:2] mux_tree_tapbuf_size5_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_30_sram;
wire [0:2] mux_tree_tapbuf_size5_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_31_sram;
wire [0:2] mux_tree_tapbuf_size5_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_32_sram;
wire [0:2] mux_tree_tapbuf_size5_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_33_sram;
wire [0:2] mux_tree_tapbuf_size5_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_34_sram;
wire [0:2] mux_tree_tapbuf_size5_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_35_sram;
wire [0:2] mux_tree_tapbuf_size5_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_36_sram;
wire [0:2] mux_tree_tapbuf_size5_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_37_sram;
wire [0:2] mux_tree_tapbuf_size5_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_38_sram;
wire [0:2] mux_tree_tapbuf_size5_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_39_sram;
wire [0:2] mux_tree_tapbuf_size5_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_40_sram;
wire [0:2] mux_tree_tapbuf_size5_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_41_sram;
wire [0:2] mux_tree_tapbuf_size5_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_42_sram;
wire [0:2] mux_tree_tapbuf_size5_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_43_sram;
wire [0:2] mux_tree_tapbuf_size5_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_44_sram;
wire [0:2] mux_tree_tapbuf_size5_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_45_sram;
wire [0:2] mux_tree_tapbuf_size5_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_46_sram;
wire [0:2] mux_tree_tapbuf_size5_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_47_sram;
wire [0:2] mux_tree_tapbuf_size5_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_48_sram;
wire [0:2] mux_tree_tapbuf_size5_48_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_49_sram;
wire [0:2] mux_tree_tapbuf_size5_49_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_50_sram;
wire [0:2] mux_tree_tapbuf_size5_50_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_51_sram;
wire [0:2] mux_tree_tapbuf_size5_51_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_52_sram;
wire [0:2] mux_tree_tapbuf_size5_52_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_53_sram;
wire [0:2] mux_tree_tapbuf_size5_53_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_54_sram;
wire [0:2] mux_tree_tapbuf_size5_54_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_55_sram;
wire [0:2] mux_tree_tapbuf_size5_55_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_56_sram;
wire [0:2] mux_tree_tapbuf_size5_56_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_57_sram;
wire [0:2] mux_tree_tapbuf_size5_57_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_58_sram;
wire [0:2] mux_tree_tapbuf_size5_58_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_59_sram;
wire [0:2] mux_tree_tapbuf_size5_59_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_60_sram;
wire [0:2] mux_tree_tapbuf_size5_60_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_61_sram;
wire [0:2] mux_tree_tapbuf_size5_61_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_62_sram;
wire [0:2] mux_tree_tapbuf_size5_62_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_63_sram;
wire [0:2] mux_tree_tapbuf_size5_63_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_64_sram;
wire [0:2] mux_tree_tapbuf_size5_64_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_65_sram;
wire [0:2] mux_tree_tapbuf_size5_65_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_66_sram;
wire [0:2] mux_tree_tapbuf_size5_66_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_67_sram;
wire [0:2] mux_tree_tapbuf_size5_67_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_68_sram;
wire [0:2] mux_tree_tapbuf_size5_68_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_69_sram;
wire [0:2] mux_tree_tapbuf_size5_69_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_70_sram;
wire [0:2] mux_tree_tapbuf_size5_70_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_71_sram;
wire [0:2] mux_tree_tapbuf_size5_71_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_72_sram;
wire [0:2] mux_tree_tapbuf_size5_72_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_73_sram;
wire [0:2] mux_tree_tapbuf_size5_73_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_74_sram;
wire [0:2] mux_tree_tapbuf_size5_74_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_75_sram;
wire [0:2] mux_tree_tapbuf_size5_75_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_76_sram;
wire [0:2] mux_tree_tapbuf_size5_76_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_77_sram;
wire [0:2] mux_tree_tapbuf_size5_77_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_78_sram;
wire [0:2] mux_tree_tapbuf_size5_78_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_79_sram;
wire [0:2] mux_tree_tapbuf_size5_79_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_80_sram;
wire [0:2] mux_tree_tapbuf_size5_80_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_81_sram;
wire [0:2] mux_tree_tapbuf_size5_81_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_82_sram;
wire [0:2] mux_tree_tapbuf_size5_82_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_83_sram;
wire [0:2] mux_tree_tapbuf_size5_83_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_84_sram;
wire [0:2] mux_tree_tapbuf_size5_84_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chanx_right_in[60];
// ----- Net sink id 1 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chanx_right_in[61];
// ----- Net sink id 1 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[150] = chanx_right_in[149];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[151] = chanx_right_in[150];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[153] = chanx_right_in[152];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[154] = chanx_right_in[153];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[155] = chanx_right_in[154];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[157] = chanx_right_in[156];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[158] = chanx_right_in[157];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[159] = chanx_right_in[158];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[161] = chanx_right_in[160];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[162] = chanx_right_in[161];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[163] = chanx_right_in[162];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[165] = chanx_right_in[164];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[166] = chanx_right_in[165];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[167] = chanx_right_in[166];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[169] = chanx_right_in[168];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[170] = chanx_right_in[169];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[171] = chanx_right_in[170];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[173] = chanx_right_in[172];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[174] = chanx_right_in[173];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[175] = chanx_right_in[174];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[132] = chanx_left_in[60];
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chanx_left_in[61];
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[150] = chanx_left_in[149];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[150];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[153] = chanx_left_in[152];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[154] = chanx_left_in[153];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[154];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[157] = chanx_left_in[156];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[158] = chanx_left_in[157];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[158];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[161] = chanx_left_in[160];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[162] = chanx_left_in[161];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[163] = chanx_left_in[162];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[165] = chanx_left_in[164];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[166] = chanx_left_in[165];
// ----- Local connection due to Wire 531 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[167] = chanx_left_in[166];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[169] = chanx_left_in[168];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[170] = chanx_left_in[169];
// ----- Local connection due to Wire 535 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[171] = chanx_left_in[170];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[173] = chanx_left_in[172];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[174] = chanx_left_in[173];
// ----- Local connection due to Wire 539 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[175] = chanx_left_in[174];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
	assign chanx_left_out[61] = chany_top_out[44];
	assign chanx_left_out[62] = chany_top_out[45];
	assign chanx_right_out[61] = chany_top_out[132];
	assign chanx_right_out[62] = chany_top_out[131];
// ----- END Local output short connections -----

	mux_tree_tapbuf_size5 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[1], chanx_right_in[7], chanx_left_in[0], chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size5 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[45], chany_top_in[90], chany_top_in[135], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size5 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[46], chany_top_in[91], chany_top_in[136], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size5 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[47], chany_top_in[92], chany_top_in[137], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size5 mux_right_track_32 (
		.in({chany_top_in[3], chany_top_in[48], chany_top_in[93], chany_top_in[138], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size5 mux_right_track_40 (
		.in({chany_top_in[4], chany_top_in[49], chany_top_in[94], chany_top_in[139], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size5 mux_right_track_48 (
		.in({chany_top_in[5], chany_top_in[50], chany_top_in[95], chany_top_in[140], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size5 mux_right_track_56 (
		.in({chany_top_in[6], chany_top_in[51], chany_top_in[96], chany_top_in[141], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size5 mux_right_track_64 (
		.in({chany_top_in[7], chany_top_in[52], chany_top_in[97], chany_top_in[142], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size5 mux_right_track_72 (
		.in({chany_top_in[8], chany_top_in[53], chany_top_in[98], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size5 mux_right_track_80 (
		.in({chany_top_in[9], chany_top_in[54], chany_top_in[99], chany_top_in[144], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size5 mux_right_track_88 (
		.in({chany_top_in[10], chany_top_in[55], chany_top_in[100], chany_top_in[145], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size5 mux_right_track_96 (
		.in({chany_top_in[11], chany_top_in[56], chany_top_in[101], chany_top_in[146], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size5 mux_right_track_104 (
		.in({chany_top_in[12], chany_top_in[57], chany_top_in[102], chany_top_in[147], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size5 mux_right_track_112 (
		.in({chany_top_in[13], chany_top_in[58], chany_top_in[103], chany_top_in[148], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size5 mux_right_track_120 (
		.in({chany_top_in[14], chany_top_in[59], chany_top_in[104], chany_top_in[149], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size5 mux_right_track_128 (
		.in({chany_top_in[15], chany_top_in[60], chany_top_in[105], chany_top_in[150], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size5 mux_right_track_136 (
		.in({chany_top_in[16], chany_top_in[61], chany_top_in[106], chany_top_in[151], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size5 mux_right_track_144 (
		.in({chany_top_in[17], chany_top_in[62], chany_top_in[107], chany_top_in[152], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size5 mux_right_track_152 (
		.in({chany_top_in[18], chany_top_in[63], chany_top_in[108], chany_top_in[153], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size5 mux_right_track_160 (
		.in({chany_top_in[19], chany_top_in[64], chany_top_in[109], chany_top_in[154], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size5 mux_right_track_168 (
		.in({chany_top_in[20], chany_top_in[65], chany_top_in[110], chany_top_in[155], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size5 mux_right_track_176 (
		.in({chany_top_in[21], chany_top_in[66], chany_top_in[111], chany_top_in[156], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size5 mux_right_track_184 (
		.in({chany_top_in[22], chany_top_in[67], chany_top_in[112], chany_top_in[157], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size5 mux_right_track_192 (
		.in({chany_top_in[23], chany_top_in[68], chany_top_in[113], chany_top_in[158], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size5 mux_right_track_200 (
		.in({chany_top_in[24], chany_top_in[69], chany_top_in[114], chany_top_in[159], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size5 mux_right_track_208 (
		.in({chany_top_in[25], chany_top_in[70], chany_top_in[115], chany_top_in[160], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size5 mux_right_track_216 (
		.in({chany_top_in[26], chany_top_in[71], chany_top_in[116], chany_top_in[161], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size5 mux_right_track_224 (
		.in({chany_top_in[27], chany_top_in[72], chany_top_in[117], chany_top_in[162], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size5 mux_right_track_232 (
		.in({chany_top_in[28], chany_top_in[73], chany_top_in[118], chany_top_in[163], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_29_sram_inv[0:2]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size5 mux_right_track_240 (
		.in({chany_top_in[29], chany_top_in[74], chany_top_in[119], chany_top_in[164], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_30_sram_inv[0:2]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size5 mux_right_track_248 (
		.in({chany_top_in[30], chany_top_in[75], chany_top_in[120], chany_top_in[165], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_31_sram_inv[0:2]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size5 mux_right_track_256 (
		.in({chany_top_in[31], chany_top_in[76], chany_top_in[121], chany_top_in[166], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_32_sram_inv[0:2]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size5 mux_right_track_264 (
		.in({chany_top_in[32], chany_top_in[77], chany_top_in[122], chany_top_in[167], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_33_sram_inv[0:2]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size5 mux_right_track_272 (
		.in({chany_top_in[33], chany_top_in[78], chany_top_in[123], chany_top_in[168], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_34_sram_inv[0:2]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size5 mux_right_track_280 (
		.in({chany_top_in[34], chany_top_in[79], chany_top_in[124], chany_top_in[169], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_35_sram_inv[0:2]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size5 mux_right_track_288 (
		.in({chany_top_in[35], chany_top_in[80], chany_top_in[125], chany_top_in[170], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_36_sram_inv[0:2]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size5 mux_right_track_296 (
		.in({chany_top_in[36], chany_top_in[81], chany_top_in[126], chany_top_in[171], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_37_sram_inv[0:2]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size5 mux_right_track_304 (
		.in({chany_top_in[37], chany_top_in[82], chany_top_in[127], chany_top_in[172], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_38_sram_inv[0:2]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size5 mux_right_track_312 (
		.in({chany_top_in[38], chany_top_in[83], chany_top_in[128], chany_top_in[173], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_39_sram_inv[0:2]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size5 mux_right_track_320 (
		.in({chany_top_in[39], chany_top_in[84], chany_top_in[129], chany_top_in[174], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_40_sram_inv[0:2]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size5 mux_right_track_328 (
		.in({chany_top_in[40], chany_top_in[85], chany_top_in[130], chany_top_in[175], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_41_sram_inv[0:2]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size5 mux_right_track_336 (
		.in({chany_top_in[41], chany_top_in[86], chany_top_in[131], chany_top_in[176], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_42_sram_inv[0:2]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size5 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[45], chany_top_in[90], chany_top_in[135], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_43_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size5 mux_left_track_33 (
		.in({chany_top_in[41], chany_top_in[86], chany_top_in[131], chany_top_in[176], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_44_sram_inv[0:2]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size5 mux_left_track_41 (
		.in({chany_top_in[40], chany_top_in[85], chany_top_in[130], chany_top_in[175], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_45_sram_inv[0:2]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size5 mux_left_track_49 (
		.in({chany_top_in[39], chany_top_in[84], chany_top_in[129], chany_top_in[174], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_46_sram_inv[0:2]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size5 mux_left_track_57 (
		.in({chany_top_in[38], chany_top_in[83], chany_top_in[128], chany_top_in[173], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_47_sram_inv[0:2]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size5 mux_left_track_65 (
		.in({chany_top_in[37], chany_top_in[82], chany_top_in[127], chany_top_in[172], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_48_sram_inv[0:2]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size5 mux_left_track_73 (
		.in({chany_top_in[36], chany_top_in[81], chany_top_in[126], chany_top_in[171], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_49_sram_inv[0:2]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size5 mux_left_track_81 (
		.in({chany_top_in[35], chany_top_in[80], chany_top_in[125], chany_top_in[170], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_50_sram_inv[0:2]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size5 mux_left_track_89 (
		.in({chany_top_in[34], chany_top_in[79], chany_top_in[124], chany_top_in[169], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_51_sram_inv[0:2]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size5 mux_left_track_97 (
		.in({chany_top_in[33], chany_top_in[78], chany_top_in[123], chany_top_in[168], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_52_sram_inv[0:2]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size5 mux_left_track_105 (
		.in({chany_top_in[32], chany_top_in[77], chany_top_in[122], chany_top_in[167], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_53_sram_inv[0:2]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size5 mux_left_track_113 (
		.in({chany_top_in[31], chany_top_in[76], chany_top_in[121], chany_top_in[166], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_54_sram_inv[0:2]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size5 mux_left_track_121 (
		.in({chany_top_in[30], chany_top_in[75], chany_top_in[120], chany_top_in[165], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_55_sram_inv[0:2]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size5 mux_left_track_129 (
		.in({chany_top_in[29], chany_top_in[74], chany_top_in[119], chany_top_in[164], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_56_sram_inv[0:2]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size5 mux_left_track_137 (
		.in({chany_top_in[28], chany_top_in[73], chany_top_in[118], chany_top_in[163], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_57_sram_inv[0:2]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size5 mux_left_track_145 (
		.in({chany_top_in[27], chany_top_in[72], chany_top_in[117], chany_top_in[162], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_58_sram_inv[0:2]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size5 mux_left_track_153 (
		.in({chany_top_in[26], chany_top_in[71], chany_top_in[116], chany_top_in[161], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_59_sram_inv[0:2]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size5 mux_left_track_161 (
		.in({chany_top_in[25], chany_top_in[70], chany_top_in[115], chany_top_in[160], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_60_sram_inv[0:2]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size5 mux_left_track_169 (
		.in({chany_top_in[24], chany_top_in[69], chany_top_in[114], chany_top_in[159], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_61_sram_inv[0:2]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size5 mux_left_track_177 (
		.in({chany_top_in[23], chany_top_in[68], chany_top_in[113], chany_top_in[158], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_62_sram_inv[0:2]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size5 mux_left_track_185 (
		.in({chany_top_in[22], chany_top_in[67], chany_top_in[112], chany_top_in[157], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_63_sram_inv[0:2]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size5 mux_left_track_193 (
		.in({chany_top_in[21], chany_top_in[66], chany_top_in[111], chany_top_in[156], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_64_sram_inv[0:2]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size5 mux_left_track_201 (
		.in({chany_top_in[20], chany_top_in[65], chany_top_in[110], chany_top_in[155], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_65_sram_inv[0:2]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size5 mux_left_track_209 (
		.in({chany_top_in[19], chany_top_in[64], chany_top_in[109], chany_top_in[154], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_66_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_66_sram_inv[0:2]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size5 mux_left_track_217 (
		.in({chany_top_in[18], chany_top_in[63], chany_top_in[108], chany_top_in[153], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_67_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_67_sram_inv[0:2]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size5 mux_left_track_225 (
		.in({chany_top_in[17], chany_top_in[62], chany_top_in[107], chany_top_in[152], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_68_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_68_sram_inv[0:2]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size5 mux_left_track_233 (
		.in({chany_top_in[16], chany_top_in[61], chany_top_in[106], chany_top_in[151], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_69_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_69_sram_inv[0:2]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size5 mux_left_track_241 (
		.in({chany_top_in[15], chany_top_in[60], chany_top_in[105], chany_top_in[150], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_70_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_70_sram_inv[0:2]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size5 mux_left_track_249 (
		.in({chany_top_in[14], chany_top_in[59], chany_top_in[104], chany_top_in[149], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_71_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_71_sram_inv[0:2]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size5 mux_left_track_257 (
		.in({chany_top_in[13], chany_top_in[58], chany_top_in[103], chany_top_in[148], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_72_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_72_sram_inv[0:2]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size5 mux_left_track_265 (
		.in({chany_top_in[12], chany_top_in[57], chany_top_in[102], chany_top_in[147], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_73_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_73_sram_inv[0:2]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size5 mux_left_track_273 (
		.in({chany_top_in[11], chany_top_in[56], chany_top_in[101], chany_top_in[146], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_74_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_74_sram_inv[0:2]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size5 mux_left_track_281 (
		.in({chany_top_in[10], chany_top_in[55], chany_top_in[100], chany_top_in[145], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_75_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_75_sram_inv[0:2]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size5 mux_left_track_289 (
		.in({chany_top_in[9], chany_top_in[54], chany_top_in[99], chany_top_in[144], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size5_76_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_76_sram_inv[0:2]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size5 mux_left_track_297 (
		.in({chany_top_in[8], chany_top_in[53], chany_top_in[98], chany_top_in[143], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_77_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_77_sram_inv[0:2]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size5 mux_left_track_305 (
		.in({chany_top_in[7], chany_top_in[52], chany_top_in[97], chany_top_in[142], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_78_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_78_sram_inv[0:2]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size5 mux_left_track_313 (
		.in({chany_top_in[6], chany_top_in[51], chany_top_in[96], chany_top_in[141], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_79_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_79_sram_inv[0:2]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size5 mux_left_track_321 (
		.in({chany_top_in[5], chany_top_in[50], chany_top_in[95], chany_top_in[140], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_80_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_80_sram_inv[0:2]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size5 mux_left_track_329 (
		.in({chany_top_in[4], chany_top_in[49], chany_top_in[94], chany_top_in[139], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_81_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_81_sram_inv[0:2]),
		.out(chanx_left_out[164]));

	mux_tree_tapbuf_size5 mux_left_track_337 (
		.in({chany_top_in[3], chany_top_in[48], chany_top_in[93], chany_top_in[138], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_82_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_82_sram_inv[0:2]),
		.out(chanx_left_out[168]));

	mux_tree_tapbuf_size5 mux_left_track_345 (
		.in({chany_top_in[2], chany_top_in[47], chany_top_in[92], chany_top_in[137], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_83_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_83_sram_inv[0:2]),
		.out(chanx_left_out[172]));

	mux_tree_tapbuf_size5 mux_left_track_353 (
		.in({chany_top_in[1], chany_top_in[46], chany_top_in[91], chany_top_in[136], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_84_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_84_sram_inv[0:2]),
		.out(chanx_left_out[176]));

	mux_tree_tapbuf_size5_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_29_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_30_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_31_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_32_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_33_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_34_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_35_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_36_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_37_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_38_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_39_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_40_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_41_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_42_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_43_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_44_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_45_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_46_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_47_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_48_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_49_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_50_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_51_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_52_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_53_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_54_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_55_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_56_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_57_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_58_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_59_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_60_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_61_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_62_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_63_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_64_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_65_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_66_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_66_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_67_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_67_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_68_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_68_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_69_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_69_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_70_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_70_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_71_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_71_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_72_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_72_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_73_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_73_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_74_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_74_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_75_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_75_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_76_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_76_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_77_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_77_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_78_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_78_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_79_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_79_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_80_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_80_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_81_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_81_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_82_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_82_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_83_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_83_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_83_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_84_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_84_sram_inv[0:2]));

	mux_tree_tapbuf_size3 mux_top_track_2 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[2], chanx_right_in[11]}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_size3 mux_top_track_38 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[26], chanx_right_in[83]}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_size3 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[28], chanx_right_in[87]}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size3 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[38], chanx_right_in[119]}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size3 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[41], chanx_right_in[127]}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_tree_tapbuf_size3 mux_top_track_74 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[50], chanx_right_in[155]}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_tree_tapbuf_size3 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[54], chanx_right_in[167]}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size3 mux_top_track_92 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[62], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chany_top_out[46]));

	mux_tree_tapbuf_size3 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[68], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chany_top_out[50]));

	mux_tree_tapbuf_size3 mux_top_track_110 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[74], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_size3 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[81], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size3 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[86], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size3 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[94], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chany_top_out[70]));

	mux_tree_tapbuf_size3 mux_top_track_146 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[98], chanx_left_in[138]}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_tree_tapbuf_size3 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[108], chanx_left_in[129]}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size3 mux_top_track_164 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[110], chanx_left_in[126]}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chany_top_out[82]));

	mux_tree_tapbuf_size3 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[121], chanx_left_in[116]}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chany_top_out[90]));

	mux_tree_tapbuf_size3 mux_top_track_182 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[122], chanx_left_in[114]}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chany_top_out[91]));

	mux_tree_tapbuf_size3 mux_top_track_218 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[146], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_top_out[109]));

	mux_tree_tapbuf_size3 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[148], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_top_out[110]));

	mux_tree_tapbuf_size3 mux_top_track_236 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[158], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_top_out[118]));

	mux_tree_tapbuf_size3 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[161], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size3 mux_top_track_254 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[170], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_top_out[127]));

	mux_tree_tapbuf_size3 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[174], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_top_out[130]));

	mux_tree_tapbuf_size3 mux_top_track_272 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[54], chanx_left_in[167]}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size3 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[49], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size3 mux_top_track_290 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[42], chanx_left_in[131]}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_top_out[145]));

	mux_tree_tapbuf_size3 mux_top_track_300 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[36], chanx_left_in[111]}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_top_out[150]));

	mux_tree_tapbuf_size3 mux_top_track_308 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[30], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_top_out[154]));

	mux_tree_tapbuf_size3 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[22], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size3 mux_top_track_326 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[18], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chany_top_out[163]));

	mux_tree_tapbuf_size3 mux_top_track_340 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[9], chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chany_top_out[170]));

	mux_tree_tapbuf_size3 mux_top_track_344 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[6], chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size3_mem mem_top_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_218 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_220 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_236 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_254 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_260 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_290 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_300 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_308 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_326 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_340 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size2 mux_top_track_4 (
		.in({chanx_right_in[4], chanx_right_in[15]}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_size2 mux_top_track_6 (
		.in({chanx_right_in[5], chanx_right_in[19]}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_size2 mux_top_track_8 (
		.in({chanx_right_in[6], chanx_right_in[23]}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size2 mux_top_track_10 (
		.in({chanx_right_in[8], chanx_right_in[27]}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_size2 mux_top_track_12 (
		.in({chanx_right_in[9], chanx_right_in[31]}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_size2 mux_top_track_14 (
		.in({chanx_right_in[10], chanx_right_in[35]}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_size2 mux_top_track_16 (
		.in({chanx_right_in[12], chanx_right_in[39]}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size2 mux_top_track_18 (
		.in({chanx_right_in[13], chanx_right_in[43]}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_size2 mux_top_track_22 (
		.in({chanx_right_in[16], chanx_right_in[51]}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_size2 mux_top_track_24 (
		.in({chanx_right_in[17], chanx_right_in[55]}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size2 mux_top_track_26 (
		.in({chanx_right_in[18], chanx_right_in[59]}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_size2 mux_top_track_28 (
		.in({chanx_right_in[20], chanx_right_in[63]}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_size2 mux_top_track_30 (
		.in({chanx_right_in[21], chanx_right_in[67]}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_size2 mux_top_track_32 (
		.in({chanx_right_in[22], chanx_right_in[71]}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size2 mux_top_track_34 (
		.in({chanx_right_in[24], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_size2 mux_top_track_36 (
		.in({chanx_right_in[25], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_size2 mux_top_track_42 (
		.in({chanx_right_in[29], chanx_right_in[91]}),
		.sram(mux_tree_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_tree_tapbuf_size2 mux_top_track_44 (
		.in({chanx_right_in[30], chanx_right_in[95]}),
		.sram(mux_tree_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_tree_tapbuf_size2 mux_top_track_46 (
		.in({chanx_right_in[32], chanx_right_in[99]}),
		.sram(mux_tree_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_18_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_size2 mux_top_track_48 (
		.in({chanx_right_in[33], chanx_right_in[103]}),
		.sram(mux_tree_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_19_sram_inv[0:1]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size2 mux_top_track_50 (
		.in({chanx_right_in[34], chanx_right_in[107]}),
		.sram(mux_tree_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_20_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_tree_tapbuf_size2 mux_top_track_52 (
		.in({chanx_right_in[36], chanx_right_in[111]}),
		.sram(mux_tree_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_21_sram_inv[0:1]),
		.out(chany_top_out[26]));

	mux_tree_tapbuf_size2 mux_top_track_54 (
		.in({chanx_right_in[37], chanx_right_in[115]}),
		.sram(mux_tree_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_22_sram_inv[0:1]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_size2 mux_top_track_58 (
		.in({chanx_right_in[40], chanx_right_in[123]}),
		.sram(mux_tree_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_23_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_tree_tapbuf_size2 mux_top_track_62 (
		.in({chanx_right_in[42], chanx_right_in[131]}),
		.sram(mux_tree_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_24_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_size2 mux_top_track_64 (
		.in({chanx_right_in[44], chanx_right_in[135]}),
		.sram(mux_tree_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_25_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size2 mux_top_track_66 (
		.in({chanx_right_in[45], chanx_right_in[139]}),
		.sram(mux_tree_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_26_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_tree_tapbuf_size2 mux_top_track_68 (
		.in({chanx_right_in[46], chanx_right_in[143]}),
		.sram(mux_tree_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_27_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_tree_tapbuf_size2 mux_top_track_70 (
		.in({chanx_right_in[48], chanx_right_in[147]}),
		.sram(mux_tree_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_28_sram_inv[0:1]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_size2 mux_top_track_72 (
		.in({chanx_right_in[49], chanx_right_in[151]}),
		.sram(mux_tree_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_29_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size2 mux_top_track_76 (
		.in({chanx_right_in[52], chanx_right_in[159]}),
		.sram(mux_tree_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_30_sram_inv[0:1]),
		.out(chany_top_out[38]));

	mux_tree_tapbuf_size2 mux_top_track_78 (
		.in({chanx_right_in[53], chanx_right_in[163]}),
		.sram(mux_tree_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_31_sram_inv[0:1]),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_size2 mux_top_track_82 (
		.in({chanx_right_in[56], chanx_right_in[171]}),
		.sram(mux_tree_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_32_sram_inv[0:1]),
		.out(chany_top_out[41]));

	mux_tree_tapbuf_size2 mux_top_track_84 (
		.in({chanx_right_in[57], chanx_right_in[175]}),
		.sram(mux_tree_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_33_sram_inv[0:1]),
		.out(chany_top_out[42]));

	mux_tree_tapbuf_size2 mux_top_track_86 (
		.in({chanx_right_in[58], chanx_right_in[176]}),
		.sram(mux_tree_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_34_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_size2 mux_top_track_94 (
		.in({chanx_right_in[64], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_35_sram_inv[0:1]),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_size2 mux_top_track_96 (
		.in({chanx_right_in[65], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_36_sram_inv[0:1]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size2 mux_top_track_98 (
		.in({chanx_right_in[66], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_37_sram_inv[0:1]),
		.out(chany_top_out[49]));

	mux_tree_tapbuf_size2 mux_top_track_102 (
		.in({chanx_right_in[69], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_38_sram_inv[0:1]),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_size2 mux_top_track_104 (
		.in({chanx_right_in[70], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_39_sram_inv[0:1]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size2 mux_top_track_106 (
		.in({chanx_right_in[72], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_40_sram_inv[0:1]),
		.out(chany_top_out[53]));

	mux_tree_tapbuf_size2 mux_top_track_108 (
		.in({chanx_right_in[73], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_41_sram_inv[0:1]),
		.out(chany_top_out[54]));

	mux_tree_tapbuf_size2 mux_top_track_112 (
		.in({chanx_right_in[76], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_42_sram_inv[0:1]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size2 mux_top_track_114 (
		.in({chanx_right_in[77], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_43_sram_inv[0:1]),
		.out(chany_top_out[57]));

	mux_tree_tapbuf_size2 mux_top_track_116 (
		.in({chanx_right_in[78], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_44_sram_inv[0:1]),
		.out(chany_top_out[58]));

	mux_tree_tapbuf_size2 mux_top_track_118 (
		.in({chanx_right_in[80], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_45_sram_inv[0:1]),
		.out(chany_top_out[59]));

	mux_tree_tapbuf_size2 mux_top_track_122 (
		.in({chanx_right_in[82], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_46_sram_inv[0:1]),
		.out(chany_top_out[61]));

	mux_tree_tapbuf_size2 mux_top_track_124 (
		.in({chanx_right_in[84], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_47_sram_inv[0:1]),
		.out(chany_top_out[62]));

	mux_tree_tapbuf_size2 mux_top_track_126 (
		.in({chanx_right_in[85], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_48_sram_inv[0:1]),
		.out(chany_top_out[63]));

	mux_tree_tapbuf_size2 mux_top_track_130 (
		.in({chanx_right_in[88], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_49_sram_inv[0:1]),
		.out(chany_top_out[65]));

	mux_tree_tapbuf_size2 mux_top_track_132 (
		.in({chanx_right_in[89], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_50_sram_inv[0:1]),
		.out(chany_top_out[66]));

	mux_tree_tapbuf_size2 mux_top_track_134 (
		.in({chanx_right_in[90], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_51_sram_inv[0:1]),
		.out(chany_top_out[67]));

	mux_tree_tapbuf_size2 mux_top_track_136 (
		.in({chanx_right_in[92], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_52_sram_inv[0:1]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size2 mux_top_track_138 (
		.in({chanx_right_in[93], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_53_sram_inv[0:1]),
		.out(chany_top_out[69]));

	mux_tree_tapbuf_size2 mux_top_track_142 (
		.in({chanx_right_in[96], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_54_sram_inv[0:1]),
		.out(chany_top_out[71]));

	mux_tree_tapbuf_size2 mux_top_track_144 (
		.in({chanx_right_in[97], chanx_left_in[140]}),
		.sram(mux_tree_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_55_sram_inv[0:1]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size2 mux_top_track_148 (
		.in({chanx_right_in[100], chanx_left_in[137]}),
		.sram(mux_tree_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_56_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_tree_tapbuf_size2 mux_top_track_150 (
		.in({chanx_right_in[101], chanx_left_in[136]}),
		.sram(mux_tree_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_57_sram_inv[0:1]),
		.out(chany_top_out[75]));

	mux_tree_tapbuf_size2 mux_top_track_152 (
		.in({chanx_right_in[102], chanx_left_in[134]}),
		.sram(mux_tree_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_58_sram_inv[0:1]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size2 mux_top_track_154 (
		.in({chanx_right_in[104], chanx_left_in[133]}),
		.sram(mux_tree_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_59_sram_inv[0:1]),
		.out(chany_top_out[77]));

	mux_tree_tapbuf_size2 mux_top_track_156 (
		.in({chanx_right_in[105], chanx_left_in[132]}),
		.sram(mux_tree_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_60_sram_inv[0:1]),
		.out(chany_top_out[78]));

	mux_tree_tapbuf_size2 mux_top_track_158 (
		.in({chanx_right_in[106], chanx_left_in[130]}),
		.sram(mux_tree_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_61_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_tree_tapbuf_size2 mux_top_track_162 (
		.in({chanx_right_in[109], chanx_left_in[128]}),
		.sram(mux_tree_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_62_sram_inv[0:1]),
		.out(chany_top_out[81]));

	mux_tree_tapbuf_size2 mux_top_track_166 (
		.in({chanx_right_in[112], chanx_left_in[125]}),
		.sram(mux_tree_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_63_sram_inv[0:1]),
		.out(chany_top_out[83]));

	mux_tree_tapbuf_size2 mux_top_track_168 (
		.in({chanx_right_in[113], chanx_left_in[124]}),
		.sram(mux_tree_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_64_sram_inv[0:1]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size2 mux_top_track_170 (
		.in({chanx_right_in[114], chanx_left_in[122]}),
		.sram(mux_tree_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_65_sram_inv[0:1]),
		.out(chany_top_out[85]));

	mux_tree_tapbuf_size2 mux_top_track_172 (
		.in({chanx_right_in[116], chanx_left_in[121]}),
		.sram(mux_tree_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_66_sram_inv[0:1]),
		.out(chany_top_out[86]));

	mux_tree_tapbuf_size2 mux_top_track_174 (
		.in({chanx_right_in[117], chanx_left_in[120]}),
		.sram(mux_tree_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_67_sram_inv[0:1]),
		.out(chany_top_out[87]));

	mux_tree_tapbuf_size2 mux_top_track_176 (
		.in({chanx_right_in[118], chanx_left_in[118]}),
		.sram(mux_tree_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_68_sram_inv[0:1]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size2 mux_top_track_178 (
		.in({chanx_right_in[120], chanx_left_in[117]}),
		.sram(mux_tree_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_69_sram_inv[0:1]),
		.out(chany_top_out[89]));

	mux_tree_tapbuf_size2 mux_top_track_184 (
		.in({chanx_right_in[124], chanx_left_in[113]}),
		.sram(mux_tree_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_70_sram_inv[0:1]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size2 mux_top_track_186 (
		.in({chanx_right_in[125], chanx_left_in[112]}),
		.sram(mux_tree_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_71_sram_inv[0:1]),
		.out(chany_top_out[93]));

	mux_tree_tapbuf_size2 mux_top_track_188 (
		.in({chanx_right_in[126], chanx_left_in[110]}),
		.sram(mux_tree_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_72_sram_inv[0:1]),
		.out(chany_top_out[94]));

	mux_tree_tapbuf_size2 mux_top_track_190 (
		.in({chanx_right_in[128], chanx_left_in[109]}),
		.sram(mux_tree_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_73_sram_inv[0:1]),
		.out(chany_top_out[95]));

	mux_tree_tapbuf_size2 mux_top_track_192 (
		.in({chanx_right_in[129], chanx_left_in[108]}),
		.sram(mux_tree_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_74_sram_inv[0:1]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size2 mux_top_track_194 (
		.in({chanx_right_in[130], chanx_left_in[106]}),
		.sram(mux_tree_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_75_sram_inv[0:1]),
		.out(chany_top_out[97]));

	mux_tree_tapbuf_size2 mux_top_track_196 (
		.in({chanx_right_in[132], chanx_left_in[105]}),
		.sram(mux_tree_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_76_sram_inv[0:1]),
		.out(chany_top_out[98]));

	mux_tree_tapbuf_size2 mux_top_track_198 (
		.in({chanx_right_in[133], chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_77_sram_inv[0:1]),
		.out(chany_top_out[99]));

	mux_tree_tapbuf_size2 mux_top_track_202 (
		.in({chanx_right_in[136], chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_78_sram_inv[0:1]),
		.out(chany_top_out[101]));

	mux_tree_tapbuf_size2 mux_top_track_204 (
		.in({chanx_right_in[137], chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_79_sram_inv[0:1]),
		.out(chany_top_out[102]));

	mux_tree_tapbuf_size2 mux_top_track_206 (
		.in({chanx_right_in[138], chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_80_sram_inv[0:1]),
		.out(chany_top_out[103]));

	mux_tree_tapbuf_size2 mux_top_track_208 (
		.in({chanx_right_in[140], chanx_left_in[97]}),
		.sram(mux_tree_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_81_sram_inv[0:1]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size2 mux_top_track_210 (
		.in({chanx_right_in[141], chanx_left_in[96]}),
		.sram(mux_tree_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_82_sram_inv[0:1]),
		.out(chany_top_out[105]));

	mux_tree_tapbuf_size2 mux_top_track_212 (
		.in({chanx_right_in[142], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_83_sram_inv[0:1]),
		.out(chany_top_out[106]));

	mux_tree_tapbuf_size2 mux_top_track_214 (
		.in({chanx_right_in[144], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_84_sram_inv[0:1]),
		.out(chany_top_out[107]));

	mux_tree_tapbuf_size2 mux_top_track_216 (
		.in({chanx_right_in[145], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_85_sram_inv[0:1]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size2 mux_top_track_222 (
		.in({chanx_right_in[149], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_86_sram_inv[0:1]),
		.out(chany_top_out[111]));

	mux_tree_tapbuf_size2 mux_top_track_224 (
		.in({chanx_right_in[150], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_87_sram_inv[0:1]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size2 mux_top_track_226 (
		.in({chanx_right_in[152], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_88_sram_inv[0:1]),
		.out(chany_top_out[113]));

	mux_tree_tapbuf_size2 mux_top_track_228 (
		.in({chanx_right_in[153], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_89_sram_inv[0:1]),
		.out(chany_top_out[114]));

	mux_tree_tapbuf_size2 mux_top_track_230 (
		.in({chanx_right_in[154], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_90_sram_inv[0:1]),
		.out(chany_top_out[115]));

	mux_tree_tapbuf_size2 mux_top_track_232 (
		.in({chanx_right_in[156], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_91_sram_inv[0:1]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size2 mux_top_track_234 (
		.in({chanx_right_in[157], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_92_sram_inv[0:1]),
		.out(chany_top_out[117]));

	mux_tree_tapbuf_size2 mux_top_track_238 (
		.in({chanx_right_in[160], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_93_sram_inv[0:1]),
		.out(chany_top_out[119]));

	mux_tree_tapbuf_size2 mux_top_track_242 (
		.in({chanx_right_in[162], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_94_sram_inv[0:1]),
		.out(chany_top_out[121]));

	mux_tree_tapbuf_size2 mux_top_track_244 (
		.in({chanx_right_in[164], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_95_sram_inv[0:1]),
		.out(chany_top_out[122]));

	mux_tree_tapbuf_size2 mux_top_track_246 (
		.in({chanx_right_in[165], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_96_sram_inv[0:1]),
		.out(chany_top_out[123]));

	mux_tree_tapbuf_size2 mux_top_track_248 (
		.in({chanx_right_in[166], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_97_sram_inv[0:1]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size2 mux_top_track_250 (
		.in({chanx_right_in[168], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_98_sram_inv[0:1]),
		.out(chany_top_out[125]));

	mux_tree_tapbuf_size2 mux_top_track_252 (
		.in({chanx_right_in[169], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_99_sram_inv[0:1]),
		.out(chany_top_out[126]));

	mux_tree_tapbuf_size2 mux_top_track_256 (
		.in({chanx_right_in[172], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_100_sram_inv[0:1]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size2 mux_top_track_258 (
		.in({chanx_right_in[173], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_101_sram_inv[0:1]),
		.out(chany_top_out[129]));

	mux_tree_tapbuf_size2 mux_top_track_266 (
		.in({chanx_left_in[58], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_102_sram_inv[0:1]),
		.out(chany_top_out[133]));

	mux_tree_tapbuf_size2 mux_top_track_268 (
		.in({chanx_left_in[57], chanx_left_in[175]}),
		.sram(mux_tree_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_103_sram_inv[0:1]),
		.out(chany_top_out[134]));

	mux_tree_tapbuf_size2 mux_top_track_270 (
		.in({chanx_left_in[56], chanx_left_in[171]}),
		.sram(mux_tree_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_104_sram_inv[0:1]),
		.out(chany_top_out[135]));

	mux_tree_tapbuf_size2 mux_top_track_274 (
		.in({chanx_left_in[53], chanx_left_in[163]}),
		.sram(mux_tree_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_105_sram_inv[0:1]),
		.out(chany_top_out[137]));

	mux_tree_tapbuf_size2 mux_top_track_276 (
		.in({chanx_left_in[52], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_106_sram_inv[0:1]),
		.out(chany_top_out[138]));

	mux_tree_tapbuf_size2 mux_top_track_278 (
		.in({chanx_left_in[50], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_107_sram_inv[0:1]),
		.out(chany_top_out[139]));

	mux_tree_tapbuf_size2 mux_top_track_282 (
		.in({chanx_left_in[48], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_108_sram_inv[0:1]),
		.out(chany_top_out[141]));

	mux_tree_tapbuf_size2 mux_top_track_284 (
		.in({chanx_left_in[46], chanx_left_in[143]}),
		.sram(mux_tree_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_109_sram_inv[0:1]),
		.out(chany_top_out[142]));

	mux_tree_tapbuf_size2 mux_top_track_286 (
		.in({chanx_left_in[45], chanx_left_in[139]}),
		.sram(mux_tree_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_110_sram_inv[0:1]),
		.out(chany_top_out[143]));

	mux_tree_tapbuf_size2 mux_top_track_288 (
		.in({chanx_left_in[44], chanx_left_in[135]}),
		.sram(mux_tree_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_111_sram_inv[0:1]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size2 mux_top_track_292 (
		.in({chanx_left_in[41], chanx_left_in[127]}),
		.sram(mux_tree_tapbuf_size2_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_112_sram_inv[0:1]),
		.out(chany_top_out[146]));

	mux_tree_tapbuf_size2 mux_top_track_294 (
		.in({chanx_left_in[40], chanx_left_in[123]}),
		.sram(mux_tree_tapbuf_size2_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_113_sram_inv[0:1]),
		.out(chany_top_out[147]));

	mux_tree_tapbuf_size2 mux_top_track_296 (
		.in({chanx_left_in[38], chanx_left_in[119]}),
		.sram(mux_tree_tapbuf_size2_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_114_sram_inv[0:1]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size2 mux_top_track_298 (
		.in({chanx_left_in[37], chanx_left_in[115]}),
		.sram(mux_tree_tapbuf_size2_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_115_sram_inv[0:1]),
		.out(chany_top_out[149]));

	mux_tree_tapbuf_size2 mux_top_track_302 (
		.in({chanx_left_in[34], chanx_left_in[107]}),
		.sram(mux_tree_tapbuf_size2_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_116_sram_inv[0:1]),
		.out(chany_top_out[151]));

	mux_tree_tapbuf_size2 mux_top_track_304 (
		.in({chanx_left_in[33], chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size2_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_117_sram_inv[0:1]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size2 mux_top_track_306 (
		.in({chanx_left_in[32], chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size2_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_118_sram_inv[0:1]),
		.out(chany_top_out[153]));

	mux_tree_tapbuf_size2 mux_top_track_310 (
		.in({chanx_left_in[29], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_size2_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_119_sram_inv[0:1]),
		.out(chany_top_out[155]));

	mux_tree_tapbuf_size2 mux_top_track_312 (
		.in({chanx_left_in[28], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_size2_120_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_120_sram_inv[0:1]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size2 mux_top_track_314 (
		.in({chanx_left_in[26], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_size2_121_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_121_sram_inv[0:1]),
		.out(chany_top_out[157]));

	mux_tree_tapbuf_size2 mux_top_track_316 (
		.in({chanx_left_in[25], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_size2_122_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_122_sram_inv[0:1]),
		.out(chany_top_out[158]));

	mux_tree_tapbuf_size2 mux_top_track_318 (
		.in({chanx_left_in[24], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_size2_123_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_123_sram_inv[0:1]),
		.out(chany_top_out[159]));

	mux_tree_tapbuf_size2 mux_top_track_322 (
		.in({chanx_left_in[21], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_size2_124_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_124_sram_inv[0:1]),
		.out(chany_top_out[161]));

	mux_tree_tapbuf_size2 mux_top_track_324 (
		.in({chanx_left_in[20], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_size2_125_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_125_sram_inv[0:1]),
		.out(chany_top_out[162]));

	mux_tree_tapbuf_size2 mux_top_track_328 (
		.in({chanx_left_in[17], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_size2_126_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_126_sram_inv[0:1]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size2 mux_top_track_330 (
		.in({chanx_left_in[16], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_size2_127_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_127_sram_inv[0:1]),
		.out(chany_top_out[165]));

	mux_tree_tapbuf_size2 mux_top_track_332 (
		.in({chanx_left_in[14], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_size2_128_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_128_sram_inv[0:1]),
		.out(chany_top_out[166]));

	mux_tree_tapbuf_size2 mux_top_track_334 (
		.in({chanx_left_in[13], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_size2_129_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_129_sram_inv[0:1]),
		.out(chany_top_out[167]));

	mux_tree_tapbuf_size2 mux_top_track_336 (
		.in({chanx_left_in[12], chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_size2_130_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_130_sram_inv[0:1]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size2 mux_top_track_338 (
		.in({chanx_left_in[10], chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_size2_131_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_131_sram_inv[0:1]),
		.out(chany_top_out[169]));

	mux_tree_tapbuf_size2 mux_top_track_342 (
		.in({chanx_left_in[8], chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_size2_132_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_132_sram_inv[0:1]),
		.out(chany_top_out[171]));

	mux_tree_tapbuf_size2 mux_top_track_346 (
		.in({chanx_left_in[5], chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_size2_133_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_133_sram_inv[0:1]),
		.out(chany_top_out[173]));

	mux_tree_tapbuf_size2 mux_top_track_348 (
		.in({chanx_left_in[4], chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_size2_134_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_134_sram_inv[0:1]),
		.out(chany_top_out[174]));

	mux_tree_tapbuf_size2 mux_top_track_350 (
		.in({chanx_left_in[2], chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_size2_135_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_135_sram_inv[0:1]),
		.out(chany_top_out[175]));

	mux_tree_tapbuf_size2_mem mem_top_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_27_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_28_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_29_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_30_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_31_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_32_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_33_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_34_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_35_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_36_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_37_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_38_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_39_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_40_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_41_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_42_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_43_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_44_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_45_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_46_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_47_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_48_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_49_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_50_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_51_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_52_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_53_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_54_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_55_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_56_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_57_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_58_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_59_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_60_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_61_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_62_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_63_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_64_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_65_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_66_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_67_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_68_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_69_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_70_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_71_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_72_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_73_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_74_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_75_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_76_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_77_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_78_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_79_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_80_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_81_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_82_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_212 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_83_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_214 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_84_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_85_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_222 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_86_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_87_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_226 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_88_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_228 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_89_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_230 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_90_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_91_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_234 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_92_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_238 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_93_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_242 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_94_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_244 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_95_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_246 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_96_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_97_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_250 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_98_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_252 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_99_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_100_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_258 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_101_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_266 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_102_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_268 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_103_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_270 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_104_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_274 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_105_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_276 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_106_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_278 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_107_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_282 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_108_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_284 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_109_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_286 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_110_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_111_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_292 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_112_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_294 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_113_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_114_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_298 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_115_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_302 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_116_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_117_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_306 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_118_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_310 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_119_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_120_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_120_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_314 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_121_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_121_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_316 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_122_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_122_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_318 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_123_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_123_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_322 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_124_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_124_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_324 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_125_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_125_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_126_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_126_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_330 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_127_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_127_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_332 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_128_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_128_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_334 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_129_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_129_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_130_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_130_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_338 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_131_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_131_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_342 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_132_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_132_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_346 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_133_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_133_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_348 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_134_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_134_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_350 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_135_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_135_sram_inv[0:1]));

	mux_tree_tapbuf_size4 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[14], chanx_right_in[47]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_size4 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[134], chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size4 mux_top_track_352 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_left_in[1], chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size4 mux_right_track_0 (
		.in({chany_top_in[44], chany_top_in[89], chany_top_in[134], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size4 mux_right_track_344 (
		.in({chany_top_in[42], chany_top_in[87], chany_top_in[132], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_4_sram_inv[0:2]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size4 mux_right_track_352 (
		.in({chany_top_in[43], chany_top_in[88], chany_top_in[133], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_5_sram_inv[0:2]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size4 mux_left_track_9 (
		.in({chany_top_in[44], chany_top_in[89], chany_top_in[134], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_6_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size4 mux_left_track_17 (
		.in({chany_top_in[43], chany_top_in[88], chany_top_in[133], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_7_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size4 mux_left_track_25 (
		.in({chany_top_in[42], chany_top_in[87], chany_top_in[132], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_8_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size4_mem mem_top_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_4_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_5_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_6_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_7_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_8_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_1__0_ -----

//----- Default net type -----
`default_nettype wire



