//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: router_bench
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Jul 24 20:28:29 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

module router_bench_top_formal_verification (
input [0:0] idata_0_0_,
input [0:0] idata_0_1_,
input [0:0] idata_0_2_,
input [0:0] idata_0_3_,
input [0:0] idata_0_4_,
input [0:0] idata_0_5_,
input [0:0] idata_0_6_,
input [0:0] idata_0_7_,
input [0:0] idata_0_8_,
input [0:0] idata_0_9_,
input [0:0] idata_0_10_,
input [0:0] idata_0_11_,
input [0:0] idata_0_12_,
input [0:0] idata_0_13_,
input [0:0] idata_0_14_,
input [0:0] idata_0_15_,
input [0:0] idata_0_16_,
input [0:0] idata_0_17_,
input [0:0] idata_0_18_,
input [0:0] idata_0_19_,
input [0:0] idata_0_20_,
input [0:0] idata_0_21_,
input [0:0] idata_0_22_,
input [0:0] idata_0_23_,
input [0:0] idata_0_24_,
input [0:0] idata_0_25_,
input [0:0] idata_0_26_,
input [0:0] idata_0_27_,
input [0:0] idata_0_28_,
input [0:0] idata_0_29_,
input [0:0] idata_0_30_,
input [0:0] idata_0_31_,
input [0:0] idata_0_32_,
input [0:0] idata_0_33_,
input [0:0] idata_0_34_,
input [0:0] ivalid_0,
input [0:0] ivch_0,
input [0:0] idata_1_0_,
input [0:0] idata_1_1_,
input [0:0] idata_1_2_,
input [0:0] idata_1_3_,
input [0:0] idata_1_4_,
input [0:0] idata_1_5_,
input [0:0] idata_1_6_,
input [0:0] idata_1_7_,
input [0:0] idata_1_8_,
input [0:0] idata_1_9_,
input [0:0] idata_1_10_,
input [0:0] idata_1_11_,
input [0:0] idata_1_12_,
input [0:0] idata_1_13_,
input [0:0] idata_1_14_,
input [0:0] idata_1_15_,
input [0:0] idata_1_16_,
input [0:0] idata_1_17_,
input [0:0] idata_1_18_,
input [0:0] idata_1_19_,
input [0:0] idata_1_20_,
input [0:0] idata_1_21_,
input [0:0] idata_1_22_,
input [0:0] idata_1_23_,
input [0:0] idata_1_24_,
input [0:0] idata_1_25_,
input [0:0] idata_1_26_,
input [0:0] idata_1_27_,
input [0:0] idata_1_28_,
input [0:0] idata_1_29_,
input [0:0] idata_1_30_,
input [0:0] idata_1_31_,
input [0:0] idata_1_32_,
input [0:0] idata_1_33_,
input [0:0] idata_1_34_,
input [0:0] ivalid_1,
input [0:0] ivch_1,
input [0:0] idata_2_0_,
input [0:0] idata_2_1_,
input [0:0] idata_2_2_,
input [0:0] idata_2_3_,
input [0:0] idata_2_4_,
input [0:0] idata_2_5_,
input [0:0] idata_2_6_,
input [0:0] idata_2_7_,
input [0:0] idata_2_8_,
input [0:0] idata_2_9_,
input [0:0] idata_2_10_,
input [0:0] idata_2_11_,
input [0:0] idata_2_12_,
input [0:0] idata_2_13_,
input [0:0] idata_2_14_,
input [0:0] idata_2_15_,
input [0:0] idata_2_16_,
input [0:0] idata_2_17_,
input [0:0] idata_2_18_,
input [0:0] idata_2_19_,
input [0:0] idata_2_20_,
input [0:0] idata_2_21_,
input [0:0] idata_2_22_,
input [0:0] idata_2_23_,
input [0:0] idata_2_24_,
input [0:0] idata_2_25_,
input [0:0] idata_2_26_,
input [0:0] idata_2_27_,
input [0:0] idata_2_28_,
input [0:0] idata_2_29_,
input [0:0] idata_2_30_,
input [0:0] idata_2_31_,
input [0:0] idata_2_32_,
input [0:0] idata_2_33_,
input [0:0] idata_2_34_,
input [0:0] ivalid_2,
input [0:0] ivch_2,
input [0:0] idata_3_0_,
input [0:0] idata_3_1_,
input [0:0] idata_3_2_,
input [0:0] idata_3_3_,
input [0:0] idata_3_4_,
input [0:0] idata_3_5_,
input [0:0] idata_3_6_,
input [0:0] idata_3_7_,
input [0:0] idata_3_8_,
input [0:0] idata_3_9_,
input [0:0] idata_3_10_,
input [0:0] idata_3_11_,
input [0:0] idata_3_12_,
input [0:0] idata_3_13_,
input [0:0] idata_3_14_,
input [0:0] idata_3_15_,
input [0:0] idata_3_16_,
input [0:0] idata_3_17_,
input [0:0] idata_3_18_,
input [0:0] idata_3_19_,
input [0:0] idata_3_20_,
input [0:0] idata_3_21_,
input [0:0] idata_3_22_,
input [0:0] idata_3_23_,
input [0:0] idata_3_24_,
input [0:0] idata_3_25_,
input [0:0] idata_3_26_,
input [0:0] idata_3_27_,
input [0:0] idata_3_28_,
input [0:0] idata_3_29_,
input [0:0] idata_3_30_,
input [0:0] idata_3_31_,
input [0:0] idata_3_32_,
input [0:0] idata_3_33_,
input [0:0] idata_3_34_,
input [0:0] ivalid_3,
input [0:0] ivch_3,
input [0:0] idata_4_0_,
input [0:0] idata_4_1_,
input [0:0] idata_4_2_,
input [0:0] idata_4_3_,
input [0:0] idata_4_4_,
input [0:0] idata_4_5_,
input [0:0] idata_4_6_,
input [0:0] idata_4_7_,
input [0:0] idata_4_8_,
input [0:0] idata_4_9_,
input [0:0] idata_4_10_,
input [0:0] idata_4_11_,
input [0:0] idata_4_12_,
input [0:0] idata_4_13_,
input [0:0] idata_4_14_,
input [0:0] idata_4_15_,
input [0:0] idata_4_16_,
input [0:0] idata_4_17_,
input [0:0] idata_4_18_,
input [0:0] idata_4_19_,
input [0:0] idata_4_20_,
input [0:0] idata_4_21_,
input [0:0] idata_4_22_,
input [0:0] idata_4_23_,
input [0:0] idata_4_24_,
input [0:0] idata_4_25_,
input [0:0] idata_4_26_,
input [0:0] idata_4_27_,
input [0:0] idata_4_28_,
input [0:0] idata_4_29_,
input [0:0] idata_4_30_,
input [0:0] idata_4_31_,
input [0:0] idata_4_32_,
input [0:0] idata_4_33_,
input [0:0] idata_4_34_,
input [0:0] ivalid_4,
input [0:0] ivch_4,
input [0:0] iack_0_0_,
input [0:0] iack_0_1_,
input [0:0] ilck_0_0_,
input [0:0] ilck_0_1_,
input [0:0] iack_1_0_,
input [0:0] iack_1_1_,
input [0:0] ilck_1_0_,
input [0:0] ilck_1_1_,
input [0:0] iack_2_0_,
input [0:0] iack_2_1_,
input [0:0] ilck_2_0_,
input [0:0] ilck_2_1_,
input [0:0] iack_3_0_,
input [0:0] iack_3_1_,
input [0:0] ilck_3_0_,
input [0:0] ilck_3_1_,
input [0:0] iack_4_0_,
input [0:0] iack_4_1_,
input [0:0] ilck_4_0_,
input [0:0] ilck_4_1_,
input [0:0] my_xpos_0_,
input [0:0] my_xpos_1_,
input [0:0] my_ypos_0_,
input [0:0] my_ypos_1_,
input [0:0] clk,
input [0:0] rst_,
output [0:0] oack_0_0_,
output [0:0] oack_0_1_,
output [0:0] ordy_0_0_,
output [0:0] ordy_0_1_,
output [0:0] olck_0_0_,
output [0:0] olck_0_1_,
output [0:0] oack_1_0_,
output [0:0] oack_1_1_,
output [0:0] ordy_1_0_,
output [0:0] ordy_1_1_,
output [0:0] olck_1_0_,
output [0:0] olck_1_1_,
output [0:0] oack_2_0_,
output [0:0] oack_2_1_,
output [0:0] ordy_2_0_,
output [0:0] ordy_2_1_,
output [0:0] olck_2_0_,
output [0:0] olck_2_1_,
output [0:0] oack_3_0_,
output [0:0] oack_3_1_,
output [0:0] ordy_3_0_,
output [0:0] ordy_3_1_,
output [0:0] olck_3_0_,
output [0:0] olck_3_1_,
output [0:0] oack_4_0_,
output [0:0] oack_4_1_,
output [0:0] ordy_4_0_,
output [0:0] ordy_4_1_,
output [0:0] olck_4_0_,
output [0:0] olck_4_1_,
output [0:0] odata_0_0_,
output [0:0] odata_0_1_,
output [0:0] odata_0_2_,
output [0:0] odata_0_3_,
output [0:0] odata_0_4_,
output [0:0] odata_0_5_,
output [0:0] odata_0_6_,
output [0:0] odata_0_7_,
output [0:0] odata_0_8_,
output [0:0] odata_0_9_,
output [0:0] odata_0_10_,
output [0:0] odata_0_11_,
output [0:0] odata_0_12_,
output [0:0] odata_0_13_,
output [0:0] odata_0_14_,
output [0:0] odata_0_15_,
output [0:0] odata_0_16_,
output [0:0] odata_0_17_,
output [0:0] odata_0_18_,
output [0:0] odata_0_19_,
output [0:0] odata_0_20_,
output [0:0] odata_0_21_,
output [0:0] odata_0_22_,
output [0:0] odata_0_23_,
output [0:0] odata_0_24_,
output [0:0] odata_0_25_,
output [0:0] odata_0_26_,
output [0:0] odata_0_27_,
output [0:0] odata_0_28_,
output [0:0] odata_0_29_,
output [0:0] odata_0_30_,
output [0:0] odata_0_31_,
output [0:0] odata_0_32_,
output [0:0] odata_0_33_,
output [0:0] odata_0_34_,
output [0:0] ovalid_0,
output [0:0] ovch_0,
output [0:0] odata_1_0_,
output [0:0] odata_1_1_,
output [0:0] odata_1_2_,
output [0:0] odata_1_3_,
output [0:0] odata_1_4_,
output [0:0] odata_1_5_,
output [0:0] odata_1_6_,
output [0:0] odata_1_7_,
output [0:0] odata_1_8_,
output [0:0] odata_1_9_,
output [0:0] odata_1_10_,
output [0:0] odata_1_11_,
output [0:0] odata_1_12_,
output [0:0] odata_1_13_,
output [0:0] odata_1_14_,
output [0:0] odata_1_15_,
output [0:0] odata_1_16_,
output [0:0] odata_1_17_,
output [0:0] odata_1_18_,
output [0:0] odata_1_19_,
output [0:0] odata_1_20_,
output [0:0] odata_1_21_,
output [0:0] odata_1_22_,
output [0:0] odata_1_23_,
output [0:0] odata_1_24_,
output [0:0] odata_1_25_,
output [0:0] odata_1_26_,
output [0:0] odata_1_27_,
output [0:0] odata_1_28_,
output [0:0] odata_1_29_,
output [0:0] odata_1_30_,
output [0:0] odata_1_31_,
output [0:0] odata_1_32_,
output [0:0] odata_1_33_,
output [0:0] odata_1_34_,
output [0:0] ovalid_1,
output [0:0] ovch_1,
output [0:0] odata_2_0_,
output [0:0] odata_2_1_,
output [0:0] odata_2_2_,
output [0:0] odata_2_3_,
output [0:0] odata_2_4_,
output [0:0] odata_2_5_,
output [0:0] odata_2_6_,
output [0:0] odata_2_7_,
output [0:0] odata_2_8_,
output [0:0] odata_2_9_,
output [0:0] odata_2_10_,
output [0:0] odata_2_11_,
output [0:0] odata_2_12_,
output [0:0] odata_2_13_,
output [0:0] odata_2_14_,
output [0:0] odata_2_15_,
output [0:0] odata_2_16_,
output [0:0] odata_2_17_,
output [0:0] odata_2_18_,
output [0:0] odata_2_19_,
output [0:0] odata_2_20_,
output [0:0] odata_2_21_,
output [0:0] odata_2_22_,
output [0:0] odata_2_23_,
output [0:0] odata_2_24_,
output [0:0] odata_2_25_,
output [0:0] odata_2_26_,
output [0:0] odata_2_27_,
output [0:0] odata_2_28_,
output [0:0] odata_2_29_,
output [0:0] odata_2_30_,
output [0:0] odata_2_31_,
output [0:0] odata_2_32_,
output [0:0] odata_2_33_,
output [0:0] odata_2_34_,
output [0:0] ovalid_2,
output [0:0] ovch_2,
output [0:0] odata_3_0_,
output [0:0] odata_3_1_,
output [0:0] odata_3_2_,
output [0:0] odata_3_3_,
output [0:0] odata_3_4_,
output [0:0] odata_3_5_,
output [0:0] odata_3_6_,
output [0:0] odata_3_7_,
output [0:0] odata_3_8_,
output [0:0] odata_3_9_,
output [0:0] odata_3_10_,
output [0:0] odata_3_11_,
output [0:0] odata_3_12_,
output [0:0] odata_3_13_,
output [0:0] odata_3_14_,
output [0:0] odata_3_15_,
output [0:0] odata_3_16_,
output [0:0] odata_3_17_,
output [0:0] odata_3_18_,
output [0:0] odata_3_19_,
output [0:0] odata_3_20_,
output [0:0] odata_3_21_,
output [0:0] odata_3_22_,
output [0:0] odata_3_23_,
output [0:0] odata_3_24_,
output [0:0] odata_3_25_,
output [0:0] odata_3_26_,
output [0:0] odata_3_27_,
output [0:0] odata_3_28_,
output [0:0] odata_3_29_,
output [0:0] odata_3_30_,
output [0:0] odata_3_31_,
output [0:0] odata_3_32_,
output [0:0] odata_3_33_,
output [0:0] odata_3_34_,
output [0:0] ovalid_3,
output [0:0] ovch_3,
output [0:0] odata_4_0_,
output [0:0] odata_4_1_,
output [0:0] odata_4_2_,
output [0:0] odata_4_3_,
output [0:0] odata_4_4_,
output [0:0] odata_4_5_,
output [0:0] odata_4_6_,
output [0:0] odata_4_7_,
output [0:0] odata_4_8_,
output [0:0] odata_4_9_,
output [0:0] odata_4_10_,
output [0:0] odata_4_11_,
output [0:0] odata_4_12_,
output [0:0] odata_4_13_,
output [0:0] odata_4_14_,
output [0:0] odata_4_15_,
output [0:0] odata_4_16_,
output [0:0] odata_4_17_,
output [0:0] odata_4_18_,
output [0:0] odata_4_19_,
output [0:0] odata_4_20_,
output [0:0] odata_4_21_,
output [0:0] odata_4_22_,
output [0:0] odata_4_23_,
output [0:0] odata_4_24_,
output [0:0] odata_4_25_,
output [0:0] odata_4_26_,
output [0:0] odata_4_27_,
output [0:0] odata_4_28_,
output [0:0] odata_4_29_,
output [0:0] odata_4_30_,
output [0:0] odata_4_31_,
output [0:0] odata_4_32_,
output [0:0] odata_4_33_,
output [0:0] odata_4_34_,
output [0:0] ovalid_4,
output [0:0] ovch_4);

// ----- Local wires for FPGA fabric -----
wire [0:479] gfpga_pad_GPIO_PAD_fm;
wire [0:0] ccff_head_fm;
wire [0:0] ccff_tail_fm;
wire [0:0] prog_clk_fm;
wire [0:0] set_fm;
wire [0:0] reset_fm;
wire [0:0] clk_fm;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		prog_clk_fm[0],
		set_fm[0],
		reset_fm[0],
		clk_fm[0],
		gfpga_pad_GPIO_PAD_fm[0:479],
		ccff_head_fm[0],
		ccff_tail_fm[0]);

// ----- Begin Connect Global ports of FPGA top module -----
	assign set_fm[0] = 1'b0;
	assign reset_fm[0] = 1'b0;
	assign clk_fm[0] = clk[0];
	assign prog_clk_fm[0] = 1'b0;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input idata_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[63] -----
	assign gfpga_pad_GPIO_PAD_fm[63] = idata_0_0_[0];

// ----- Blif Benchmark input idata_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[88] -----
	assign gfpga_pad_GPIO_PAD_fm[88] = idata_0_1_[0];

// ----- Blif Benchmark input idata_0_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[467] -----
	assign gfpga_pad_GPIO_PAD_fm[467] = idata_0_2_[0];

// ----- Blif Benchmark input idata_0_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[162] -----
	assign gfpga_pad_GPIO_PAD_fm[162] = idata_0_3_[0];

// ----- Blif Benchmark input idata_0_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[303] -----
	assign gfpga_pad_GPIO_PAD_fm[303] = idata_0_4_[0];

// ----- Blif Benchmark input idata_0_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[67] -----
	assign gfpga_pad_GPIO_PAD_fm[67] = idata_0_5_[0];

// ----- Blif Benchmark input idata_0_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[167] -----
	assign gfpga_pad_GPIO_PAD_fm[167] = idata_0_6_[0];

// ----- Blif Benchmark input idata_0_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[463] -----
	assign gfpga_pad_GPIO_PAD_fm[463] = idata_0_7_[0];

// ----- Blif Benchmark input idata_0_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[106] -----
	assign gfpga_pad_GPIO_PAD_fm[106] = idata_0_8_[0];

// ----- Blif Benchmark input idata_0_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[182] -----
	assign gfpga_pad_GPIO_PAD_fm[182] = idata_0_9_[0];

// ----- Blif Benchmark input idata_0_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[71] -----
	assign gfpga_pad_GPIO_PAD_fm[71] = idata_0_10_[0];

// ----- Blif Benchmark input idata_0_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[33] -----
	assign gfpga_pad_GPIO_PAD_fm[33] = idata_0_11_[0];

// ----- Blif Benchmark input idata_0_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[195] -----
	assign gfpga_pad_GPIO_PAD_fm[195] = idata_0_12_[0];

// ----- Blif Benchmark input idata_0_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[310] -----
	assign gfpga_pad_GPIO_PAD_fm[310] = idata_0_13_[0];

// ----- Blif Benchmark input idata_0_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[29] -----
	assign gfpga_pad_GPIO_PAD_fm[29] = idata_0_14_[0];

// ----- Blif Benchmark input idata_0_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[331] -----
	assign gfpga_pad_GPIO_PAD_fm[331] = idata_0_15_[0];

// ----- Blif Benchmark input idata_0_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[356] -----
	assign gfpga_pad_GPIO_PAD_fm[356] = idata_0_16_[0];

// ----- Blif Benchmark input idata_0_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[249] -----
	assign gfpga_pad_GPIO_PAD_fm[249] = idata_0_17_[0];

// ----- Blif Benchmark input idata_0_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[289] -----
	assign gfpga_pad_GPIO_PAD_fm[289] = idata_0_18_[0];

// ----- Blif Benchmark input idata_0_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[418] -----
	assign gfpga_pad_GPIO_PAD_fm[418] = idata_0_19_[0];

// ----- Blif Benchmark input idata_0_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[436] -----
	assign gfpga_pad_GPIO_PAD_fm[436] = idata_0_20_[0];

// ----- Blif Benchmark input idata_0_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[387] -----
	assign gfpga_pad_GPIO_PAD_fm[387] = idata_0_21_[0];

// ----- Blif Benchmark input idata_0_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[60] -----
	assign gfpga_pad_GPIO_PAD_fm[60] = idata_0_22_[0];

// ----- Blif Benchmark input idata_0_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[361] -----
	assign gfpga_pad_GPIO_PAD_fm[361] = idata_0_23_[0];

// ----- Blif Benchmark input idata_0_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[231] -----
	assign gfpga_pad_GPIO_PAD_fm[231] = idata_0_24_[0];

// ----- Blif Benchmark input idata_0_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[253] -----
	assign gfpga_pad_GPIO_PAD_fm[253] = idata_0_25_[0];

// ----- Blif Benchmark input idata_0_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[252] -----
	assign gfpga_pad_GPIO_PAD_fm[252] = idata_0_26_[0];

// ----- Blif Benchmark input idata_0_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[28] -----
	assign gfpga_pad_GPIO_PAD_fm[28] = idata_0_27_[0];

// ----- Blif Benchmark input idata_0_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[408] -----
	assign gfpga_pad_GPIO_PAD_fm[408] = idata_0_28_[0];

// ----- Blif Benchmark input idata_0_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[450] -----
	assign gfpga_pad_GPIO_PAD_fm[450] = idata_0_29_[0];

// ----- Blif Benchmark input idata_0_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[178] -----
	assign gfpga_pad_GPIO_PAD_fm[178] = idata_0_30_[0];

// ----- Blif Benchmark input idata_0_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[44] -----
	assign gfpga_pad_GPIO_PAD_fm[44] = idata_0_31_[0];

// ----- Blif Benchmark input idata_0_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[455] -----
	assign gfpga_pad_GPIO_PAD_fm[455] = idata_0_32_[0];

// ----- Blif Benchmark input idata_0_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[42] -----
	assign gfpga_pad_GPIO_PAD_fm[42] = idata_0_33_[0];

// ----- Blif Benchmark input idata_0_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[40] -----
	assign gfpga_pad_GPIO_PAD_fm[40] = idata_0_34_[0];

// ----- Blif Benchmark input ivalid_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[132] -----
	assign gfpga_pad_GPIO_PAD_fm[132] = ivalid_0[0];

// ----- Blif Benchmark input ivch_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[388] -----
	assign gfpga_pad_GPIO_PAD_fm[388] = ivch_0[0];

// ----- Blif Benchmark input idata_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[327] -----
	assign gfpga_pad_GPIO_PAD_fm[327] = idata_1_0_[0];

// ----- Blif Benchmark input idata_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[55] -----
	assign gfpga_pad_GPIO_PAD_fm[55] = idata_1_1_[0];

// ----- Blif Benchmark input idata_1_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[176] -----
	assign gfpga_pad_GPIO_PAD_fm[176] = idata_1_2_[0];

// ----- Blif Benchmark input idata_1_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[120] -----
	assign gfpga_pad_GPIO_PAD_fm[120] = idata_1_3_[0];

// ----- Blif Benchmark input idata_1_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[272] -----
	assign gfpga_pad_GPIO_PAD_fm[272] = idata_1_4_[0];

// ----- Blif Benchmark input idata_1_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[30] -----
	assign gfpga_pad_GPIO_PAD_fm[30] = idata_1_5_[0];

// ----- Blif Benchmark input idata_1_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[473] -----
	assign gfpga_pad_GPIO_PAD_fm[473] = idata_1_6_[0];

// ----- Blif Benchmark input idata_1_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[59] -----
	assign gfpga_pad_GPIO_PAD_fm[59] = idata_1_7_[0];

// ----- Blif Benchmark input idata_1_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[232] -----
	assign gfpga_pad_GPIO_PAD_fm[232] = idata_1_8_[0];

// ----- Blif Benchmark input idata_1_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[448] -----
	assign gfpga_pad_GPIO_PAD_fm[448] = idata_1_9_[0];

// ----- Blif Benchmark input idata_1_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[370] -----
	assign gfpga_pad_GPIO_PAD_fm[370] = idata_1_10_[0];

// ----- Blif Benchmark input idata_1_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[111] -----
	assign gfpga_pad_GPIO_PAD_fm[111] = idata_1_11_[0];

// ----- Blif Benchmark input idata_1_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[292] -----
	assign gfpga_pad_GPIO_PAD_fm[292] = idata_1_12_[0];

// ----- Blif Benchmark input idata_1_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[144] -----
	assign gfpga_pad_GPIO_PAD_fm[144] = idata_1_13_[0];

// ----- Blif Benchmark input idata_1_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[209] -----
	assign gfpga_pad_GPIO_PAD_fm[209] = idata_1_14_[0];

// ----- Blif Benchmark input idata_1_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[61] -----
	assign gfpga_pad_GPIO_PAD_fm[61] = idata_1_15_[0];

// ----- Blif Benchmark input idata_1_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[13] -----
	assign gfpga_pad_GPIO_PAD_fm[13] = idata_1_16_[0];

// ----- Blif Benchmark input idata_1_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[27] -----
	assign gfpga_pad_GPIO_PAD_fm[27] = idata_1_17_[0];

// ----- Blif Benchmark input idata_1_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[228] -----
	assign gfpga_pad_GPIO_PAD_fm[228] = idata_1_18_[0];

// ----- Blif Benchmark input idata_1_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[288] -----
	assign gfpga_pad_GPIO_PAD_fm[288] = idata_1_19_[0];

// ----- Blif Benchmark input idata_1_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[194] -----
	assign gfpga_pad_GPIO_PAD_fm[194] = idata_1_20_[0];

// ----- Blif Benchmark input idata_1_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[18] -----
	assign gfpga_pad_GPIO_PAD_fm[18] = idata_1_21_[0];

// ----- Blif Benchmark input idata_1_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[131] -----
	assign gfpga_pad_GPIO_PAD_fm[131] = idata_1_22_[0];

// ----- Blif Benchmark input idata_1_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[449] -----
	assign gfpga_pad_GPIO_PAD_fm[449] = idata_1_23_[0];

// ----- Blif Benchmark input idata_1_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[113] -----
	assign gfpga_pad_GPIO_PAD_fm[113] = idata_1_24_[0];

// ----- Blif Benchmark input idata_1_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[165] -----
	assign gfpga_pad_GPIO_PAD_fm[165] = idata_1_25_[0];

// ----- Blif Benchmark input idata_1_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[333] -----
	assign gfpga_pad_GPIO_PAD_fm[333] = idata_1_26_[0];

// ----- Blif Benchmark input idata_1_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[406] -----
	assign gfpga_pad_GPIO_PAD_fm[406] = idata_1_27_[0];

// ----- Blif Benchmark input idata_1_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[3] -----
	assign gfpga_pad_GPIO_PAD_fm[3] = idata_1_28_[0];

// ----- Blif Benchmark input idata_1_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[35] -----
	assign gfpga_pad_GPIO_PAD_fm[35] = idata_1_29_[0];

// ----- Blif Benchmark input idata_1_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[200] -----
	assign gfpga_pad_GPIO_PAD_fm[200] = idata_1_30_[0];

// ----- Blif Benchmark input idata_1_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[280] -----
	assign gfpga_pad_GPIO_PAD_fm[280] = idata_1_31_[0];

// ----- Blif Benchmark input idata_1_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[365] -----
	assign gfpga_pad_GPIO_PAD_fm[365] = idata_1_32_[0];

// ----- Blif Benchmark input idata_1_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[420] -----
	assign gfpga_pad_GPIO_PAD_fm[420] = idata_1_33_[0];

// ----- Blif Benchmark input idata_1_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[335] -----
	assign gfpga_pad_GPIO_PAD_fm[335] = idata_1_34_[0];

// ----- Blif Benchmark input ivalid_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[97] -----
	assign gfpga_pad_GPIO_PAD_fm[97] = ivalid_1[0];

// ----- Blif Benchmark input ivch_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[32] -----
	assign gfpga_pad_GPIO_PAD_fm[32] = ivch_1[0];

// ----- Blif Benchmark input idata_2_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[142] -----
	assign gfpga_pad_GPIO_PAD_fm[142] = idata_2_0_[0];

// ----- Blif Benchmark input idata_2_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[155] -----
	assign gfpga_pad_GPIO_PAD_fm[155] = idata_2_1_[0];

// ----- Blif Benchmark input idata_2_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[99] -----
	assign gfpga_pad_GPIO_PAD_fm[99] = idata_2_2_[0];

// ----- Blif Benchmark input idata_2_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[39] -----
	assign gfpga_pad_GPIO_PAD_fm[39] = idata_2_3_[0];

// ----- Blif Benchmark input idata_2_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[238] -----
	assign gfpga_pad_GPIO_PAD_fm[238] = idata_2_4_[0];

// ----- Blif Benchmark input idata_2_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[326] -----
	assign gfpga_pad_GPIO_PAD_fm[326] = idata_2_5_[0];

// ----- Blif Benchmark input idata_2_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[186] -----
	assign gfpga_pad_GPIO_PAD_fm[186] = idata_2_6_[0];

// ----- Blif Benchmark input idata_2_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[187] -----
	assign gfpga_pad_GPIO_PAD_fm[187] = idata_2_7_[0];

// ----- Blif Benchmark input idata_2_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[123] -----
	assign gfpga_pad_GPIO_PAD_fm[123] = idata_2_8_[0];

// ----- Blif Benchmark input idata_2_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[402] -----
	assign gfpga_pad_GPIO_PAD_fm[402] = idata_2_9_[0];

// ----- Blif Benchmark input idata_2_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[193] -----
	assign gfpga_pad_GPIO_PAD_fm[193] = idata_2_10_[0];

// ----- Blif Benchmark input idata_2_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[429] -----
	assign gfpga_pad_GPIO_PAD_fm[429] = idata_2_11_[0];

// ----- Blif Benchmark input idata_2_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[282] -----
	assign gfpga_pad_GPIO_PAD_fm[282] = idata_2_12_[0];

// ----- Blif Benchmark input idata_2_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[304] -----
	assign gfpga_pad_GPIO_PAD_fm[304] = idata_2_13_[0];

// ----- Blif Benchmark input idata_2_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[283] -----
	assign gfpga_pad_GPIO_PAD_fm[283] = idata_2_14_[0];

// ----- Blif Benchmark input idata_2_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[206] -----
	assign gfpga_pad_GPIO_PAD_fm[206] = idata_2_15_[0];

// ----- Blif Benchmark input idata_2_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[295] -----
	assign gfpga_pad_GPIO_PAD_fm[295] = idata_2_16_[0];

// ----- Blif Benchmark input idata_2_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[366] -----
	assign gfpga_pad_GPIO_PAD_fm[366] = idata_2_17_[0];

// ----- Blif Benchmark input idata_2_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[259] -----
	assign gfpga_pad_GPIO_PAD_fm[259] = idata_2_18_[0];

// ----- Blif Benchmark input idata_2_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[457] -----
	assign gfpga_pad_GPIO_PAD_fm[457] = idata_2_19_[0];

// ----- Blif Benchmark input idata_2_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[362] -----
	assign gfpga_pad_GPIO_PAD_fm[362] = idata_2_20_[0];

// ----- Blif Benchmark input idata_2_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[469] -----
	assign gfpga_pad_GPIO_PAD_fm[469] = idata_2_21_[0];

// ----- Blif Benchmark input idata_2_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[125] -----
	assign gfpga_pad_GPIO_PAD_fm[125] = idata_2_22_[0];

// ----- Blif Benchmark input idata_2_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[390] -----
	assign gfpga_pad_GPIO_PAD_fm[390] = idata_2_23_[0];

// ----- Blif Benchmark input idata_2_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[399] -----
	assign gfpga_pad_GPIO_PAD_fm[399] = idata_2_24_[0];

// ----- Blif Benchmark input idata_2_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[299] -----
	assign gfpga_pad_GPIO_PAD_fm[299] = idata_2_25_[0];

// ----- Blif Benchmark input idata_2_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[46] -----
	assign gfpga_pad_GPIO_PAD_fm[46] = idata_2_26_[0];

// ----- Blif Benchmark input idata_2_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[81] -----
	assign gfpga_pad_GPIO_PAD_fm[81] = idata_2_27_[0];

// ----- Blif Benchmark input idata_2_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[108] -----
	assign gfpga_pad_GPIO_PAD_fm[108] = idata_2_28_[0];

// ----- Blif Benchmark input idata_2_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[379] -----
	assign gfpga_pad_GPIO_PAD_fm[379] = idata_2_29_[0];

// ----- Blif Benchmark input idata_2_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[64] -----
	assign gfpga_pad_GPIO_PAD_fm[64] = idata_2_30_[0];

// ----- Blif Benchmark input idata_2_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[373] -----
	assign gfpga_pad_GPIO_PAD_fm[373] = idata_2_31_[0];

// ----- Blif Benchmark input idata_2_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[425] -----
	assign gfpga_pad_GPIO_PAD_fm[425] = idata_2_32_[0];

// ----- Blif Benchmark input idata_2_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[135] -----
	assign gfpga_pad_GPIO_PAD_fm[135] = idata_2_33_[0];

// ----- Blif Benchmark input idata_2_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[24] -----
	assign gfpga_pad_GPIO_PAD_fm[24] = idata_2_34_[0];

// ----- Blif Benchmark input ivalid_2 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[101] -----
	assign gfpga_pad_GPIO_PAD_fm[101] = ivalid_2[0];

// ----- Blif Benchmark input ivch_2 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[409] -----
	assign gfpga_pad_GPIO_PAD_fm[409] = ivch_2[0];

// ----- Blif Benchmark input idata_3_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[296] -----
	assign gfpga_pad_GPIO_PAD_fm[296] = idata_3_0_[0];

// ----- Blif Benchmark input idata_3_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[460] -----
	assign gfpga_pad_GPIO_PAD_fm[460] = idata_3_1_[0];

// ----- Blif Benchmark input idata_3_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[31] -----
	assign gfpga_pad_GPIO_PAD_fm[31] = idata_3_2_[0];

// ----- Blif Benchmark input idata_3_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[103] -----
	assign gfpga_pad_GPIO_PAD_fm[103] = idata_3_3_[0];

// ----- Blif Benchmark input idata_3_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[277] -----
	assign gfpga_pad_GPIO_PAD_fm[277] = idata_3_4_[0];

// ----- Blif Benchmark input idata_3_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[382] -----
	assign gfpga_pad_GPIO_PAD_fm[382] = idata_3_5_[0];

// ----- Blif Benchmark input idata_3_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[404] -----
	assign gfpga_pad_GPIO_PAD_fm[404] = idata_3_6_[0];

// ----- Blif Benchmark input idata_3_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[171] -----
	assign gfpga_pad_GPIO_PAD_fm[171] = idata_3_7_[0];

// ----- Blif Benchmark input idata_3_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[281] -----
	assign gfpga_pad_GPIO_PAD_fm[281] = idata_3_8_[0];

// ----- Blif Benchmark input idata_3_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[349] -----
	assign gfpga_pad_GPIO_PAD_fm[349] = idata_3_9_[0];

// ----- Blif Benchmark input idata_3_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[439] -----
	assign gfpga_pad_GPIO_PAD_fm[439] = idata_3_10_[0];

// ----- Blif Benchmark input idata_3_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[413] -----
	assign gfpga_pad_GPIO_PAD_fm[413] = idata_3_11_[0];

// ----- Blif Benchmark input idata_3_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[377] -----
	assign gfpga_pad_GPIO_PAD_fm[377] = idata_3_12_[0];

// ----- Blif Benchmark input idata_3_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[87] -----
	assign gfpga_pad_GPIO_PAD_fm[87] = idata_3_13_[0];

// ----- Blif Benchmark input idata_3_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[217] -----
	assign gfpga_pad_GPIO_PAD_fm[217] = idata_3_14_[0];

// ----- Blif Benchmark input idata_3_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[57] -----
	assign gfpga_pad_GPIO_PAD_fm[57] = idata_3_15_[0];

// ----- Blif Benchmark input idata_3_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[279] -----
	assign gfpga_pad_GPIO_PAD_fm[279] = idata_3_16_[0];

// ----- Blif Benchmark input idata_3_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[116] -----
	assign gfpga_pad_GPIO_PAD_fm[116] = idata_3_17_[0];

// ----- Blif Benchmark input idata_3_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[2] -----
	assign gfpga_pad_GPIO_PAD_fm[2] = idata_3_18_[0];

// ----- Blif Benchmark input idata_3_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[419] -----
	assign gfpga_pad_GPIO_PAD_fm[419] = idata_3_19_[0];

// ----- Blif Benchmark input idata_3_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[66] -----
	assign gfpga_pad_GPIO_PAD_fm[66] = idata_3_20_[0];

// ----- Blif Benchmark input idata_3_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[215] -----
	assign gfpga_pad_GPIO_PAD_fm[215] = idata_3_21_[0];

// ----- Blif Benchmark input idata_3_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[318] -----
	assign gfpga_pad_GPIO_PAD_fm[318] = idata_3_22_[0];

// ----- Blif Benchmark input idata_3_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[329] -----
	assign gfpga_pad_GPIO_PAD_fm[329] = idata_3_23_[0];

// ----- Blif Benchmark input idata_3_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[286] -----
	assign gfpga_pad_GPIO_PAD_fm[286] = idata_3_24_[0];

// ----- Blif Benchmark input idata_3_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[363] -----
	assign gfpga_pad_GPIO_PAD_fm[363] = idata_3_25_[0];

// ----- Blif Benchmark input idata_3_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[308] -----
	assign gfpga_pad_GPIO_PAD_fm[308] = idata_3_26_[0];

// ----- Blif Benchmark input idata_3_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[434] -----
	assign gfpga_pad_GPIO_PAD_fm[434] = idata_3_27_[0];

// ----- Blif Benchmark input idata_3_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[173] -----
	assign gfpga_pad_GPIO_PAD_fm[173] = idata_3_28_[0];

// ----- Blif Benchmark input idata_3_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[287] -----
	assign gfpga_pad_GPIO_PAD_fm[287] = idata_3_29_[0];

// ----- Blif Benchmark input idata_3_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[83] -----
	assign gfpga_pad_GPIO_PAD_fm[83] = idata_3_30_[0];

// ----- Blif Benchmark input idata_3_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[146] -----
	assign gfpga_pad_GPIO_PAD_fm[146] = idata_3_31_[0];

// ----- Blif Benchmark input idata_3_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[328] -----
	assign gfpga_pad_GPIO_PAD_fm[328] = idata_3_32_[0];

// ----- Blif Benchmark input idata_3_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[380] -----
	assign gfpga_pad_GPIO_PAD_fm[380] = idata_3_33_[0];

// ----- Blif Benchmark input idata_3_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[17] -----
	assign gfpga_pad_GPIO_PAD_fm[17] = idata_3_34_[0];

// ----- Blif Benchmark input ivalid_3 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[74] -----
	assign gfpga_pad_GPIO_PAD_fm[74] = ivalid_3[0];

// ----- Blif Benchmark input ivch_3 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[414] -----
	assign gfpga_pad_GPIO_PAD_fm[414] = ivch_3[0];

// ----- Blif Benchmark input idata_4_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[133] -----
	assign gfpga_pad_GPIO_PAD_fm[133] = idata_4_0_[0];

// ----- Blif Benchmark input idata_4_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[112] -----
	assign gfpga_pad_GPIO_PAD_fm[112] = idata_4_1_[0];

// ----- Blif Benchmark input idata_4_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[300] -----
	assign gfpga_pad_GPIO_PAD_fm[300] = idata_4_2_[0];

// ----- Blif Benchmark input idata_4_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[188] -----
	assign gfpga_pad_GPIO_PAD_fm[188] = idata_4_3_[0];

// ----- Blif Benchmark input idata_4_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[265] -----
	assign gfpga_pad_GPIO_PAD_fm[265] = idata_4_4_[0];

// ----- Blif Benchmark input idata_4_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[130] -----
	assign gfpga_pad_GPIO_PAD_fm[130] = idata_4_5_[0];

// ----- Blif Benchmark input idata_4_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[38] -----
	assign gfpga_pad_GPIO_PAD_fm[38] = idata_4_6_[0];

// ----- Blif Benchmark input idata_4_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[158] -----
	assign gfpga_pad_GPIO_PAD_fm[158] = idata_4_7_[0];

// ----- Blif Benchmark input idata_4_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[451] -----
	assign gfpga_pad_GPIO_PAD_fm[451] = idata_4_8_[0];

// ----- Blif Benchmark input idata_4_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[405] -----
	assign gfpga_pad_GPIO_PAD_fm[405] = idata_4_9_[0];

// ----- Blif Benchmark input idata_4_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[201] -----
	assign gfpga_pad_GPIO_PAD_fm[201] = idata_4_10_[0];

// ----- Blif Benchmark input idata_4_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[92] -----
	assign gfpga_pad_GPIO_PAD_fm[92] = idata_4_11_[0];

// ----- Blif Benchmark input idata_4_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[179] -----
	assign gfpga_pad_GPIO_PAD_fm[179] = idata_4_12_[0];

// ----- Blif Benchmark input idata_4_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[266] -----
	assign gfpga_pad_GPIO_PAD_fm[266] = idata_4_13_[0];

// ----- Blif Benchmark input idata_4_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[431] -----
	assign gfpga_pad_GPIO_PAD_fm[431] = idata_4_14_[0];

// ----- Blif Benchmark input idata_4_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[4] -----
	assign gfpga_pad_GPIO_PAD_fm[4] = idata_4_15_[0];

// ----- Blif Benchmark input idata_4_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[330] -----
	assign gfpga_pad_GPIO_PAD_fm[330] = idata_4_16_[0];

// ----- Blif Benchmark input idata_4_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[474] -----
	assign gfpga_pad_GPIO_PAD_fm[474] = idata_4_17_[0];

// ----- Blif Benchmark input idata_4_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[203] -----
	assign gfpga_pad_GPIO_PAD_fm[203] = idata_4_18_[0];

// ----- Blif Benchmark input idata_4_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[397] -----
	assign gfpga_pad_GPIO_PAD_fm[397] = idata_4_19_[0];

// ----- Blif Benchmark input idata_4_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[16] -----
	assign gfpga_pad_GPIO_PAD_fm[16] = idata_4_20_[0];

// ----- Blif Benchmark input idata_4_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[157] -----
	assign gfpga_pad_GPIO_PAD_fm[157] = idata_4_21_[0];

// ----- Blif Benchmark input idata_4_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[230] -----
	assign gfpga_pad_GPIO_PAD_fm[230] = idata_4_22_[0];

// ----- Blif Benchmark input idata_4_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[351] -----
	assign gfpga_pad_GPIO_PAD_fm[351] = idata_4_23_[0];

// ----- Blif Benchmark input idata_4_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[20] -----
	assign gfpga_pad_GPIO_PAD_fm[20] = idata_4_24_[0];

// ----- Blif Benchmark input idata_4_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[341] -----
	assign gfpga_pad_GPIO_PAD_fm[341] = idata_4_25_[0];

// ----- Blif Benchmark input idata_4_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[435] -----
	assign gfpga_pad_GPIO_PAD_fm[435] = idata_4_26_[0];

// ----- Blif Benchmark input idata_4_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[378] -----
	assign gfpga_pad_GPIO_PAD_fm[378] = idata_4_27_[0];

// ----- Blif Benchmark input idata_4_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[86] -----
	assign gfpga_pad_GPIO_PAD_fm[86] = idata_4_28_[0];

// ----- Blif Benchmark input idata_4_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[442] -----
	assign gfpga_pad_GPIO_PAD_fm[442] = idata_4_29_[0];

// ----- Blif Benchmark input idata_4_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[23] -----
	assign gfpga_pad_GPIO_PAD_fm[23] = idata_4_30_[0];

// ----- Blif Benchmark input idata_4_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[294] -----
	assign gfpga_pad_GPIO_PAD_fm[294] = idata_4_31_[0];

// ----- Blif Benchmark input idata_4_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[441] -----
	assign gfpga_pad_GPIO_PAD_fm[441] = idata_4_32_[0];

// ----- Blif Benchmark input idata_4_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[427] -----
	assign gfpga_pad_GPIO_PAD_fm[427] = idata_4_33_[0];

// ----- Blif Benchmark input idata_4_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[69] -----
	assign gfpga_pad_GPIO_PAD_fm[69] = idata_4_34_[0];

// ----- Blif Benchmark input ivalid_4 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[6] -----
	assign gfpga_pad_GPIO_PAD_fm[6] = ivalid_4[0];

// ----- Blif Benchmark input ivch_4 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[102] -----
	assign gfpga_pad_GPIO_PAD_fm[102] = ivch_4[0];

// ----- Blif Benchmark input iack_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[21] -----
	assign gfpga_pad_GPIO_PAD_fm[21] = iack_0_0_[0];

// ----- Blif Benchmark input iack_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[180] -----
	assign gfpga_pad_GPIO_PAD_fm[180] = iack_0_1_[0];

// ----- Blif Benchmark input ilck_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[309] -----
	assign gfpga_pad_GPIO_PAD_fm[309] = ilck_0_0_[0];

// ----- Blif Benchmark input ilck_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[411] -----
	assign gfpga_pad_GPIO_PAD_fm[411] = ilck_0_1_[0];

// ----- Blif Benchmark input iack_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[458] -----
	assign gfpga_pad_GPIO_PAD_fm[458] = iack_1_0_[0];

// ----- Blif Benchmark input iack_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[336] -----
	assign gfpga_pad_GPIO_PAD_fm[336] = iack_1_1_[0];

// ----- Blif Benchmark input ilck_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[394] -----
	assign gfpga_pad_GPIO_PAD_fm[394] = ilck_1_0_[0];

// ----- Blif Benchmark input ilck_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[352] -----
	assign gfpga_pad_GPIO_PAD_fm[352] = ilck_1_1_[0];

// ----- Blif Benchmark input iack_2_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[346] -----
	assign gfpga_pad_GPIO_PAD_fm[346] = iack_2_0_[0];

// ----- Blif Benchmark input iack_2_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[306] -----
	assign gfpga_pad_GPIO_PAD_fm[306] = iack_2_1_[0];

// ----- Blif Benchmark input ilck_2_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[79] -----
	assign gfpga_pad_GPIO_PAD_fm[79] = ilck_2_0_[0];

// ----- Blif Benchmark input ilck_2_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[219] -----
	assign gfpga_pad_GPIO_PAD_fm[219] = ilck_2_1_[0];

// ----- Blif Benchmark input iack_3_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[430] -----
	assign gfpga_pad_GPIO_PAD_fm[430] = iack_3_0_[0];

// ----- Blif Benchmark input iack_3_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[470] -----
	assign gfpga_pad_GPIO_PAD_fm[470] = iack_3_1_[0];

// ----- Blif Benchmark input ilck_3_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[267] -----
	assign gfpga_pad_GPIO_PAD_fm[267] = ilck_3_0_[0];

// ----- Blif Benchmark input ilck_3_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[53] -----
	assign gfpga_pad_GPIO_PAD_fm[53] = ilck_3_1_[0];

// ----- Blif Benchmark input iack_4_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[192] -----
	assign gfpga_pad_GPIO_PAD_fm[192] = iack_4_0_[0];

// ----- Blif Benchmark input iack_4_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[54] -----
	assign gfpga_pad_GPIO_PAD_fm[54] = iack_4_1_[0];

// ----- Blif Benchmark input ilck_4_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[177] -----
	assign gfpga_pad_GPIO_PAD_fm[177] = ilck_4_0_[0];

// ----- Blif Benchmark input ilck_4_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[396] -----
	assign gfpga_pad_GPIO_PAD_fm[396] = ilck_4_1_[0];

// ----- Blif Benchmark input my_xpos_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[340] -----
	assign gfpga_pad_GPIO_PAD_fm[340] = my_xpos_0_[0];

// ----- Blif Benchmark input my_xpos_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[143] -----
	assign gfpga_pad_GPIO_PAD_fm[143] = my_xpos_1_[0];

// ----- Blif Benchmark input my_ypos_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[159] -----
	assign gfpga_pad_GPIO_PAD_fm[159] = my_ypos_0_[0];

// ----- Blif Benchmark input my_ypos_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[8] -----
	assign gfpga_pad_GPIO_PAD_fm[8] = my_ypos_1_[0];

// ----- Blif Benchmark input clk is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[236] -----
	assign gfpga_pad_GPIO_PAD_fm[236] = clk[0];

// ----- Blif Benchmark input rst_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[211] -----
	assign gfpga_pad_GPIO_PAD_fm[211] = rst_[0];

// ----- Blif Benchmark output oack_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[41] -----
	assign oack_0_0_[0] = gfpga_pad_GPIO_PAD_fm[41];

// ----- Blif Benchmark output oack_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[14] -----
	assign oack_0_1_[0] = gfpga_pad_GPIO_PAD_fm[14];

// ----- Blif Benchmark output ordy_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[73] -----
	assign ordy_0_0_[0] = gfpga_pad_GPIO_PAD_fm[73];

// ----- Blif Benchmark output ordy_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[410] -----
	assign ordy_0_1_[0] = gfpga_pad_GPIO_PAD_fm[410];

// ----- Blif Benchmark output olck_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[472] -----
	assign olck_0_0_[0] = gfpga_pad_GPIO_PAD_fm[472];

// ----- Blif Benchmark output olck_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[244] -----
	assign olck_0_1_[0] = gfpga_pad_GPIO_PAD_fm[244];

// ----- Blif Benchmark output oack_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[478] -----
	assign oack_1_0_[0] = gfpga_pad_GPIO_PAD_fm[478];

// ----- Blif Benchmark output oack_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[354] -----
	assign oack_1_1_[0] = gfpga_pad_GPIO_PAD_fm[354];

// ----- Blif Benchmark output ordy_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[10] -----
	assign ordy_1_0_[0] = gfpga_pad_GPIO_PAD_fm[10];

// ----- Blif Benchmark output ordy_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[446] -----
	assign ordy_1_1_[0] = gfpga_pad_GPIO_PAD_fm[446];

// ----- Blif Benchmark output olck_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[461] -----
	assign olck_1_0_[0] = gfpga_pad_GPIO_PAD_fm[461];

// ----- Blif Benchmark output olck_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[109] -----
	assign olck_1_1_[0] = gfpga_pad_GPIO_PAD_fm[109];

// ----- Blif Benchmark output oack_2_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[220] -----
	assign oack_2_0_[0] = gfpga_pad_GPIO_PAD_fm[220];

// ----- Blif Benchmark output oack_2_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[437] -----
	assign oack_2_1_[0] = gfpga_pad_GPIO_PAD_fm[437];

// ----- Blif Benchmark output ordy_2_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[170] -----
	assign ordy_2_0_[0] = gfpga_pad_GPIO_PAD_fm[170];

// ----- Blif Benchmark output ordy_2_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[400] -----
	assign ordy_2_1_[0] = gfpga_pad_GPIO_PAD_fm[400];

// ----- Blif Benchmark output olck_2_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[118] -----
	assign olck_2_0_[0] = gfpga_pad_GPIO_PAD_fm[118];

// ----- Blif Benchmark output olck_2_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[70] -----
	assign olck_2_1_[0] = gfpga_pad_GPIO_PAD_fm[70];

// ----- Blif Benchmark output oack_3_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[258] -----
	assign oack_3_0_[0] = gfpga_pad_GPIO_PAD_fm[258];

// ----- Blif Benchmark output oack_3_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[138] -----
	assign oack_3_1_[0] = gfpga_pad_GPIO_PAD_fm[138];

// ----- Blif Benchmark output ordy_3_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[48] -----
	assign ordy_3_0_[0] = gfpga_pad_GPIO_PAD_fm[48];

// ----- Blif Benchmark output ordy_3_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[117] -----
	assign ordy_3_1_[0] = gfpga_pad_GPIO_PAD_fm[117];

// ----- Blif Benchmark output olck_3_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[364] -----
	assign olck_3_0_[0] = gfpga_pad_GPIO_PAD_fm[364];

// ----- Blif Benchmark output olck_3_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[190] -----
	assign olck_3_1_[0] = gfpga_pad_GPIO_PAD_fm[190];

// ----- Blif Benchmark output oack_4_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[290] -----
	assign oack_4_0_[0] = gfpga_pad_GPIO_PAD_fm[290];

// ----- Blif Benchmark output oack_4_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[381] -----
	assign oack_4_1_[0] = gfpga_pad_GPIO_PAD_fm[381];

// ----- Blif Benchmark output ordy_4_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[126] -----
	assign ordy_4_0_[0] = gfpga_pad_GPIO_PAD_fm[126];

// ----- Blif Benchmark output ordy_4_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[386] -----
	assign ordy_4_1_[0] = gfpga_pad_GPIO_PAD_fm[386];

// ----- Blif Benchmark output olck_4_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[421] -----
	assign olck_4_0_[0] = gfpga_pad_GPIO_PAD_fm[421];

// ----- Blif Benchmark output olck_4_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[104] -----
	assign olck_4_1_[0] = gfpga_pad_GPIO_PAD_fm[104];

// ----- Blif Benchmark output odata_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[127] -----
	assign odata_0_0_[0] = gfpga_pad_GPIO_PAD_fm[127];

// ----- Blif Benchmark output odata_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[82] -----
	assign odata_0_1_[0] = gfpga_pad_GPIO_PAD_fm[82];

// ----- Blif Benchmark output odata_0_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[93] -----
	assign odata_0_2_[0] = gfpga_pad_GPIO_PAD_fm[93];

// ----- Blif Benchmark output odata_0_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[302] -----
	assign odata_0_3_[0] = gfpga_pad_GPIO_PAD_fm[302];

// ----- Blif Benchmark output odata_0_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[338] -----
	assign odata_0_4_[0] = gfpga_pad_GPIO_PAD_fm[338];

// ----- Blif Benchmark output odata_0_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[260] -----
	assign odata_0_5_[0] = gfpga_pad_GPIO_PAD_fm[260];

// ----- Blif Benchmark output odata_0_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[45] -----
	assign odata_0_6_[0] = gfpga_pad_GPIO_PAD_fm[45];

// ----- Blif Benchmark output odata_0_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[12] -----
	assign odata_0_7_[0] = gfpga_pad_GPIO_PAD_fm[12];

// ----- Blif Benchmark output odata_0_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[367] -----
	assign odata_0_8_[0] = gfpga_pad_GPIO_PAD_fm[367];

// ----- Blif Benchmark output odata_0_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[212] -----
	assign odata_0_9_[0] = gfpga_pad_GPIO_PAD_fm[212];

// ----- Blif Benchmark output odata_0_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[189] -----
	assign odata_0_10_[0] = gfpga_pad_GPIO_PAD_fm[189];

// ----- Blif Benchmark output odata_0_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[447] -----
	assign odata_0_11_[0] = gfpga_pad_GPIO_PAD_fm[447];

// ----- Blif Benchmark output odata_0_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[428] -----
	assign odata_0_12_[0] = gfpga_pad_GPIO_PAD_fm[428];

// ----- Blif Benchmark output odata_0_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[174] -----
	assign odata_0_13_[0] = gfpga_pad_GPIO_PAD_fm[174];

// ----- Blif Benchmark output odata_0_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[37] -----
	assign odata_0_14_[0] = gfpga_pad_GPIO_PAD_fm[37];

// ----- Blif Benchmark output odata_0_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[114] -----
	assign odata_0_15_[0] = gfpga_pad_GPIO_PAD_fm[114];

// ----- Blif Benchmark output odata_0_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[264] -----
	assign odata_0_16_[0] = gfpga_pad_GPIO_PAD_fm[264];

// ----- Blif Benchmark output odata_0_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[293] -----
	assign odata_0_17_[0] = gfpga_pad_GPIO_PAD_fm[293];

// ----- Blif Benchmark output odata_0_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[94] -----
	assign odata_0_18_[0] = gfpga_pad_GPIO_PAD_fm[94];

// ----- Blif Benchmark output odata_0_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[355] -----
	assign odata_0_19_[0] = gfpga_pad_GPIO_PAD_fm[355];

// ----- Blif Benchmark output odata_0_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[213] -----
	assign odata_0_20_[0] = gfpga_pad_GPIO_PAD_fm[213];

// ----- Blif Benchmark output odata_0_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[433] -----
	assign odata_0_21_[0] = gfpga_pad_GPIO_PAD_fm[433];

// ----- Blif Benchmark output odata_0_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[141] -----
	assign odata_0_22_[0] = gfpga_pad_GPIO_PAD_fm[141];

// ----- Blif Benchmark output odata_0_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[43] -----
	assign odata_0_23_[0] = gfpga_pad_GPIO_PAD_fm[43];

// ----- Blif Benchmark output odata_0_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[75] -----
	assign odata_0_24_[0] = gfpga_pad_GPIO_PAD_fm[75];

// ----- Blif Benchmark output odata_0_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[274] -----
	assign odata_0_25_[0] = gfpga_pad_GPIO_PAD_fm[274];

// ----- Blif Benchmark output odata_0_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[169] -----
	assign odata_0_26_[0] = gfpga_pad_GPIO_PAD_fm[169];

// ----- Blif Benchmark output odata_0_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[185] -----
	assign odata_0_27_[0] = gfpga_pad_GPIO_PAD_fm[185];

// ----- Blif Benchmark output odata_0_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[175] -----
	assign odata_0_28_[0] = gfpga_pad_GPIO_PAD_fm[175];

// ----- Blif Benchmark output odata_0_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[369] -----
	assign odata_0_29_[0] = gfpga_pad_GPIO_PAD_fm[369];

// ----- Blif Benchmark output odata_0_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[353] -----
	assign odata_0_30_[0] = gfpga_pad_GPIO_PAD_fm[353];

// ----- Blif Benchmark output odata_0_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[214] -----
	assign odata_0_31_[0] = gfpga_pad_GPIO_PAD_fm[214];

// ----- Blif Benchmark output odata_0_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[273] -----
	assign odata_0_32_[0] = gfpga_pad_GPIO_PAD_fm[273];

// ----- Blif Benchmark output odata_0_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[471] -----
	assign odata_0_33_[0] = gfpga_pad_GPIO_PAD_fm[471];

// ----- Blif Benchmark output odata_0_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[246] -----
	assign odata_0_34_[0] = gfpga_pad_GPIO_PAD_fm[246];

// ----- Blif Benchmark output ovalid_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[383] -----
	assign ovalid_0[0] = gfpga_pad_GPIO_PAD_fm[383];

// ----- Blif Benchmark output ovch_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[395] -----
	assign ovch_0[0] = gfpga_pad_GPIO_PAD_fm[395];

// ----- Blif Benchmark output odata_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[98] -----
	assign odata_1_0_[0] = gfpga_pad_GPIO_PAD_fm[98];

// ----- Blif Benchmark output odata_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[269] -----
	assign odata_1_1_[0] = gfpga_pad_GPIO_PAD_fm[269];

// ----- Blif Benchmark output odata_1_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[15] -----
	assign odata_1_2_[0] = gfpga_pad_GPIO_PAD_fm[15];

// ----- Blif Benchmark output odata_1_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[339] -----
	assign odata_1_3_[0] = gfpga_pad_GPIO_PAD_fm[339];

// ----- Blif Benchmark output odata_1_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[107] -----
	assign odata_1_4_[0] = gfpga_pad_GPIO_PAD_fm[107];

// ----- Blif Benchmark output odata_1_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[301] -----
	assign odata_1_5_[0] = gfpga_pad_GPIO_PAD_fm[301];

// ----- Blif Benchmark output odata_1_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[342] -----
	assign odata_1_6_[0] = gfpga_pad_GPIO_PAD_fm[342];

// ----- Blif Benchmark output odata_1_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[368] -----
	assign odata_1_7_[0] = gfpga_pad_GPIO_PAD_fm[368];

// ----- Blif Benchmark output odata_1_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[77] -----
	assign odata_1_8_[0] = gfpga_pad_GPIO_PAD_fm[77];

// ----- Blif Benchmark output odata_1_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[423] -----
	assign odata_1_9_[0] = gfpga_pad_GPIO_PAD_fm[423];

// ----- Blif Benchmark output odata_1_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[191] -----
	assign odata_1_10_[0] = gfpga_pad_GPIO_PAD_fm[191];

// ----- Blif Benchmark output odata_1_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[210] -----
	assign odata_1_11_[0] = gfpga_pad_GPIO_PAD_fm[210];

// ----- Blif Benchmark output odata_1_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[459] -----
	assign odata_1_12_[0] = gfpga_pad_GPIO_PAD_fm[459];

// ----- Blif Benchmark output odata_1_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[374] -----
	assign odata_1_13_[0] = gfpga_pad_GPIO_PAD_fm[374];

// ----- Blif Benchmark output odata_1_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[137] -----
	assign odata_1_14_[0] = gfpga_pad_GPIO_PAD_fm[137];

// ----- Blif Benchmark output odata_1_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[51] -----
	assign odata_1_15_[0] = gfpga_pad_GPIO_PAD_fm[51];

// ----- Blif Benchmark output odata_1_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[348] -----
	assign odata_1_16_[0] = gfpga_pad_GPIO_PAD_fm[348];

// ----- Blif Benchmark output odata_1_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[0] -----
	assign odata_1_17_[0] = gfpga_pad_GPIO_PAD_fm[0];

// ----- Blif Benchmark output odata_1_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[65] -----
	assign odata_1_18_[0] = gfpga_pad_GPIO_PAD_fm[65];

// ----- Blif Benchmark output odata_1_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[371] -----
	assign odata_1_19_[0] = gfpga_pad_GPIO_PAD_fm[371];

// ----- Blif Benchmark output odata_1_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[168] -----
	assign odata_1_20_[0] = gfpga_pad_GPIO_PAD_fm[168];

// ----- Blif Benchmark output odata_1_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[438] -----
	assign odata_1_21_[0] = gfpga_pad_GPIO_PAD_fm[438];

// ----- Blif Benchmark output odata_1_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[1] -----
	assign odata_1_22_[0] = gfpga_pad_GPIO_PAD_fm[1];

// ----- Blif Benchmark output odata_1_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[462] -----
	assign odata_1_23_[0] = gfpga_pad_GPIO_PAD_fm[462];

// ----- Blif Benchmark output odata_1_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[26] -----
	assign odata_1_24_[0] = gfpga_pad_GPIO_PAD_fm[26];

// ----- Blif Benchmark output odata_1_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[122] -----
	assign odata_1_25_[0] = gfpga_pad_GPIO_PAD_fm[122];

// ----- Blif Benchmark output odata_1_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[372] -----
	assign odata_1_26_[0] = gfpga_pad_GPIO_PAD_fm[372];

// ----- Blif Benchmark output odata_1_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[432] -----
	assign odata_1_27_[0] = gfpga_pad_GPIO_PAD_fm[432];

// ----- Blif Benchmark output odata_1_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[464] -----
	assign odata_1_28_[0] = gfpga_pad_GPIO_PAD_fm[464];

// ----- Blif Benchmark output odata_1_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[233] -----
	assign odata_1_29_[0] = gfpga_pad_GPIO_PAD_fm[233];

// ----- Blif Benchmark output odata_1_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[222] -----
	assign odata_1_30_[0] = gfpga_pad_GPIO_PAD_fm[222];

// ----- Blif Benchmark output odata_1_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[307] -----
	assign odata_1_31_[0] = gfpga_pad_GPIO_PAD_fm[307];

// ----- Blif Benchmark output odata_1_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[344] -----
	assign odata_1_32_[0] = gfpga_pad_GPIO_PAD_fm[344];

// ----- Blif Benchmark output odata_1_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[89] -----
	assign odata_1_33_[0] = gfpga_pad_GPIO_PAD_fm[89];

// ----- Blif Benchmark output odata_1_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[454] -----
	assign odata_1_34_[0] = gfpga_pad_GPIO_PAD_fm[454];

// ----- Blif Benchmark output ovalid_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[407] -----
	assign ovalid_1[0] = gfpga_pad_GPIO_PAD_fm[407];

// ----- Blif Benchmark output ovch_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[128] -----
	assign ovch_1[0] = gfpga_pad_GPIO_PAD_fm[128];

// ----- Blif Benchmark output odata_2_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[49] -----
	assign odata_2_0_[0] = gfpga_pad_GPIO_PAD_fm[49];

// ----- Blif Benchmark output odata_2_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[322] -----
	assign odata_2_1_[0] = gfpga_pad_GPIO_PAD_fm[322];

// ----- Blif Benchmark output odata_2_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[466] -----
	assign odata_2_2_[0] = gfpga_pad_GPIO_PAD_fm[466];

// ----- Blif Benchmark output odata_2_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[199] -----
	assign odata_2_3_[0] = gfpga_pad_GPIO_PAD_fm[199];

// ----- Blif Benchmark output odata_2_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[204] -----
	assign odata_2_4_[0] = gfpga_pad_GPIO_PAD_fm[204];

// ----- Blif Benchmark output odata_2_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[181] -----
	assign odata_2_5_[0] = gfpga_pad_GPIO_PAD_fm[181];

// ----- Blif Benchmark output odata_2_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[350] -----
	assign odata_2_6_[0] = gfpga_pad_GPIO_PAD_fm[350];

// ----- Blif Benchmark output odata_2_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[166] -----
	assign odata_2_7_[0] = gfpga_pad_GPIO_PAD_fm[166];

// ----- Blif Benchmark output odata_2_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[477] -----
	assign odata_2_8_[0] = gfpga_pad_GPIO_PAD_fm[477];

// ----- Blif Benchmark output odata_2_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[62] -----
	assign odata_2_9_[0] = gfpga_pad_GPIO_PAD_fm[62];

// ----- Blif Benchmark output odata_2_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[7] -----
	assign odata_2_10_[0] = gfpga_pad_GPIO_PAD_fm[7];

// ----- Blif Benchmark output odata_2_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[453] -----
	assign odata_2_11_[0] = gfpga_pad_GPIO_PAD_fm[453];

// ----- Blif Benchmark output odata_2_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[284] -----
	assign odata_2_12_[0] = gfpga_pad_GPIO_PAD_fm[284];

// ----- Blif Benchmark output odata_2_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[25] -----
	assign odata_2_13_[0] = gfpga_pad_GPIO_PAD_fm[25];

// ----- Blif Benchmark output odata_2_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[56] -----
	assign odata_2_14_[0] = gfpga_pad_GPIO_PAD_fm[56];

// ----- Blif Benchmark output odata_2_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[268] -----
	assign odata_2_15_[0] = gfpga_pad_GPIO_PAD_fm[268];

// ----- Blif Benchmark output odata_2_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[401] -----
	assign odata_2_16_[0] = gfpga_pad_GPIO_PAD_fm[401];

// ----- Blif Benchmark output odata_2_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[129] -----
	assign odata_2_17_[0] = gfpga_pad_GPIO_PAD_fm[129];

// ----- Blif Benchmark output odata_2_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[140] -----
	assign odata_2_18_[0] = gfpga_pad_GPIO_PAD_fm[140];

// ----- Blif Benchmark output odata_2_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[263] -----
	assign odata_2_19_[0] = gfpga_pad_GPIO_PAD_fm[263];

// ----- Blif Benchmark output odata_2_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[202] -----
	assign odata_2_20_[0] = gfpga_pad_GPIO_PAD_fm[202];

// ----- Blif Benchmark output odata_2_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[391] -----
	assign odata_2_21_[0] = gfpga_pad_GPIO_PAD_fm[391];

// ----- Blif Benchmark output odata_2_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[417] -----
	assign odata_2_22_[0] = gfpga_pad_GPIO_PAD_fm[417];

// ----- Blif Benchmark output odata_2_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[50] -----
	assign odata_2_23_[0] = gfpga_pad_GPIO_PAD_fm[50];

// ----- Blif Benchmark output odata_2_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[216] -----
	assign odata_2_24_[0] = gfpga_pad_GPIO_PAD_fm[216];

// ----- Blif Benchmark output odata_2_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[312] -----
	assign odata_2_25_[0] = gfpga_pad_GPIO_PAD_fm[312];

// ----- Blif Benchmark output odata_2_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[121] -----
	assign odata_2_26_[0] = gfpga_pad_GPIO_PAD_fm[121];

// ----- Blif Benchmark output odata_2_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[343] -----
	assign odata_2_27_[0] = gfpga_pad_GPIO_PAD_fm[343];

// ----- Blif Benchmark output odata_2_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[229] -----
	assign odata_2_28_[0] = gfpga_pad_GPIO_PAD_fm[229];

// ----- Blif Benchmark output odata_2_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[139] -----
	assign odata_2_29_[0] = gfpga_pad_GPIO_PAD_fm[139];

// ----- Blif Benchmark output odata_2_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[163] -----
	assign odata_2_30_[0] = gfpga_pad_GPIO_PAD_fm[163];

// ----- Blif Benchmark output odata_2_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[151] -----
	assign odata_2_31_[0] = gfpga_pad_GPIO_PAD_fm[151];

// ----- Blif Benchmark output odata_2_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[468] -----
	assign odata_2_32_[0] = gfpga_pad_GPIO_PAD_fm[468];

// ----- Blif Benchmark output odata_2_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[398] -----
	assign odata_2_33_[0] = gfpga_pad_GPIO_PAD_fm[398];

// ----- Blif Benchmark output odata_2_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[297] -----
	assign odata_2_34_[0] = gfpga_pad_GPIO_PAD_fm[297];

// ----- Blif Benchmark output ovalid_2 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[426] -----
	assign ovalid_2[0] = gfpga_pad_GPIO_PAD_fm[426];

// ----- Blif Benchmark output ovch_2 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[376] -----
	assign ovch_2[0] = gfpga_pad_GPIO_PAD_fm[376];

// ----- Blif Benchmark output odata_3_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[403] -----
	assign odata_3_0_[0] = gfpga_pad_GPIO_PAD_fm[403];

// ----- Blif Benchmark output odata_3_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[208] -----
	assign odata_3_1_[0] = gfpga_pad_GPIO_PAD_fm[208];

// ----- Blif Benchmark output odata_3_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[218] -----
	assign odata_3_2_[0] = gfpga_pad_GPIO_PAD_fm[218];

// ----- Blif Benchmark output odata_3_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[440] -----
	assign odata_3_3_[0] = gfpga_pad_GPIO_PAD_fm[440];

// ----- Blif Benchmark output odata_3_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[19] -----
	assign odata_3_4_[0] = gfpga_pad_GPIO_PAD_fm[19];

// ----- Blif Benchmark output odata_3_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[456] -----
	assign odata_3_5_[0] = gfpga_pad_GPIO_PAD_fm[456];

// ----- Blif Benchmark output odata_3_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[58] -----
	assign odata_3_6_[0] = gfpga_pad_GPIO_PAD_fm[58];

// ----- Blif Benchmark output odata_3_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[36] -----
	assign odata_3_7_[0] = gfpga_pad_GPIO_PAD_fm[36];

// ----- Blif Benchmark output odata_3_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[124] -----
	assign odata_3_8_[0] = gfpga_pad_GPIO_PAD_fm[124];

// ----- Blif Benchmark output odata_3_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[298] -----
	assign odata_3_9_[0] = gfpga_pad_GPIO_PAD_fm[298];

// ----- Blif Benchmark output odata_3_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[11] -----
	assign odata_3_10_[0] = gfpga_pad_GPIO_PAD_fm[11];

// ----- Blif Benchmark output odata_3_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[68] -----
	assign odata_3_11_[0] = gfpga_pad_GPIO_PAD_fm[68];

// ----- Blif Benchmark output odata_3_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[337] -----
	assign odata_3_12_[0] = gfpga_pad_GPIO_PAD_fm[337];

// ----- Blif Benchmark output odata_3_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[270] -----
	assign odata_3_13_[0] = gfpga_pad_GPIO_PAD_fm[270];

// ----- Blif Benchmark output odata_3_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[285] -----
	assign odata_3_14_[0] = gfpga_pad_GPIO_PAD_fm[285];

// ----- Blif Benchmark output odata_3_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[345] -----
	assign odata_3_15_[0] = gfpga_pad_GPIO_PAD_fm[345];

// ----- Blif Benchmark output odata_3_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[9] -----
	assign odata_3_16_[0] = gfpga_pad_GPIO_PAD_fm[9];

// ----- Blif Benchmark output odata_3_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[465] -----
	assign odata_3_17_[0] = gfpga_pad_GPIO_PAD_fm[465];

// ----- Blif Benchmark output odata_3_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[452] -----
	assign odata_3_18_[0] = gfpga_pad_GPIO_PAD_fm[452];

// ----- Blif Benchmark output odata_3_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[305] -----
	assign odata_3_19_[0] = gfpga_pad_GPIO_PAD_fm[305];

// ----- Blif Benchmark output odata_3_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[254] -----
	assign odata_3_20_[0] = gfpga_pad_GPIO_PAD_fm[254];

// ----- Blif Benchmark output odata_3_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[145] -----
	assign odata_3_21_[0] = gfpga_pad_GPIO_PAD_fm[145];

// ----- Blif Benchmark output odata_3_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[445] -----
	assign odata_3_22_[0] = gfpga_pad_GPIO_PAD_fm[445];

// ----- Blif Benchmark output odata_3_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[223] -----
	assign odata_3_23_[0] = gfpga_pad_GPIO_PAD_fm[223];

// ----- Blif Benchmark output odata_3_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[52] -----
	assign odata_3_24_[0] = gfpga_pad_GPIO_PAD_fm[52];

// ----- Blif Benchmark output odata_3_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[197] -----
	assign odata_3_25_[0] = gfpga_pad_GPIO_PAD_fm[197];

// ----- Blif Benchmark output odata_3_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[196] -----
	assign odata_3_26_[0] = gfpga_pad_GPIO_PAD_fm[196];

// ----- Blif Benchmark output odata_3_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[183] -----
	assign odata_3_27_[0] = gfpga_pad_GPIO_PAD_fm[183];

// ----- Blif Benchmark output odata_3_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[291] -----
	assign odata_3_28_[0] = gfpga_pad_GPIO_PAD_fm[291];

// ----- Blif Benchmark output odata_3_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[358] -----
	assign odata_3_29_[0] = gfpga_pad_GPIO_PAD_fm[358];

// ----- Blif Benchmark output odata_3_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[422] -----
	assign odata_3_30_[0] = gfpga_pad_GPIO_PAD_fm[422];

// ----- Blif Benchmark output odata_3_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[424] -----
	assign odata_3_31_[0] = gfpga_pad_GPIO_PAD_fm[424];

// ----- Blif Benchmark output odata_3_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[476] -----
	assign odata_3_32_[0] = gfpga_pad_GPIO_PAD_fm[476];

// ----- Blif Benchmark output odata_3_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[95] -----
	assign odata_3_33_[0] = gfpga_pad_GPIO_PAD_fm[95];

// ----- Blif Benchmark output odata_3_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[359] -----
	assign odata_3_34_[0] = gfpga_pad_GPIO_PAD_fm[359];

// ----- Blif Benchmark output ovalid_3 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[221] -----
	assign ovalid_3[0] = gfpga_pad_GPIO_PAD_fm[221];

// ----- Blif Benchmark output ovch_3 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[161] -----
	assign ovch_3[0] = gfpga_pad_GPIO_PAD_fm[161];

// ----- Blif Benchmark output odata_4_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[198] -----
	assign odata_4_0_[0] = gfpga_pad_GPIO_PAD_fm[198];

// ----- Blif Benchmark output odata_4_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[393] -----
	assign odata_4_1_[0] = gfpga_pad_GPIO_PAD_fm[393];

// ----- Blif Benchmark output odata_4_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[134] -----
	assign odata_4_2_[0] = gfpga_pad_GPIO_PAD_fm[134];

// ----- Blif Benchmark output odata_4_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[392] -----
	assign odata_4_3_[0] = gfpga_pad_GPIO_PAD_fm[392];

// ----- Blif Benchmark output odata_4_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[360] -----
	assign odata_4_4_[0] = gfpga_pad_GPIO_PAD_fm[360];

// ----- Blif Benchmark output odata_4_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[385] -----
	assign odata_4_5_[0] = gfpga_pad_GPIO_PAD_fm[385];

// ----- Blif Benchmark output odata_4_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[389] -----
	assign odata_4_6_[0] = gfpga_pad_GPIO_PAD_fm[389];

// ----- Blif Benchmark output odata_4_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[416] -----
	assign odata_4_7_[0] = gfpga_pad_GPIO_PAD_fm[416];

// ----- Blif Benchmark output odata_4_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[479] -----
	assign odata_4_8_[0] = gfpga_pad_GPIO_PAD_fm[479];

// ----- Blif Benchmark output odata_4_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[275] -----
	assign odata_4_9_[0] = gfpga_pad_GPIO_PAD_fm[275];

// ----- Blif Benchmark output odata_4_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[321] -----
	assign odata_4_10_[0] = gfpga_pad_GPIO_PAD_fm[321];

// ----- Blif Benchmark output odata_4_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[100] -----
	assign odata_4_11_[0] = gfpga_pad_GPIO_PAD_fm[100];

// ----- Blif Benchmark output odata_4_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[313] -----
	assign odata_4_12_[0] = gfpga_pad_GPIO_PAD_fm[313];

// ----- Blif Benchmark output odata_4_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[34] -----
	assign odata_4_13_[0] = gfpga_pad_GPIO_PAD_fm[34];

// ----- Blif Benchmark output odata_4_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[323] -----
	assign odata_4_14_[0] = gfpga_pad_GPIO_PAD_fm[323];

// ----- Blif Benchmark output odata_4_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[207] -----
	assign odata_4_15_[0] = gfpga_pad_GPIO_PAD_fm[207];

// ----- Blif Benchmark output odata_4_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[119] -----
	assign odata_4_16_[0] = gfpga_pad_GPIO_PAD_fm[119];

// ----- Blif Benchmark output odata_4_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[72] -----
	assign odata_4_17_[0] = gfpga_pad_GPIO_PAD_fm[72];

// ----- Blif Benchmark output odata_4_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[78] -----
	assign odata_4_18_[0] = gfpga_pad_GPIO_PAD_fm[78];

// ----- Blif Benchmark output odata_4_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[110] -----
	assign odata_4_19_[0] = gfpga_pad_GPIO_PAD_fm[110];

// ----- Blif Benchmark output odata_4_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[384] -----
	assign odata_4_20_[0] = gfpga_pad_GPIO_PAD_fm[384];

// ----- Blif Benchmark output odata_4_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[105] -----
	assign odata_4_21_[0] = gfpga_pad_GPIO_PAD_fm[105];

// ----- Blif Benchmark output odata_4_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[47] -----
	assign odata_4_22_[0] = gfpga_pad_GPIO_PAD_fm[47];

// ----- Blif Benchmark output odata_4_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[115] -----
	assign odata_4_23_[0] = gfpga_pad_GPIO_PAD_fm[115];

// ----- Blif Benchmark output odata_4_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[475] -----
	assign odata_4_24_[0] = gfpga_pad_GPIO_PAD_fm[475];

// ----- Blif Benchmark output odata_4_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[357] -----
	assign odata_4_25_[0] = gfpga_pad_GPIO_PAD_fm[357];

// ----- Blif Benchmark output odata_4_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[443] -----
	assign odata_4_26_[0] = gfpga_pad_GPIO_PAD_fm[443];

// ----- Blif Benchmark output odata_4_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[271] -----
	assign odata_4_27_[0] = gfpga_pad_GPIO_PAD_fm[271];

// ----- Blif Benchmark output odata_4_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[278] -----
	assign odata_4_28_[0] = gfpga_pad_GPIO_PAD_fm[278];

// ----- Blif Benchmark output odata_4_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[160] -----
	assign odata_4_29_[0] = gfpga_pad_GPIO_PAD_fm[160];

// ----- Blif Benchmark output odata_4_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[205] -----
	assign odata_4_30_[0] = gfpga_pad_GPIO_PAD_fm[205];

// ----- Blif Benchmark output odata_4_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[136] -----
	assign odata_4_31_[0] = gfpga_pad_GPIO_PAD_fm[136];

// ----- Blif Benchmark output odata_4_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[184] -----
	assign odata_4_32_[0] = gfpga_pad_GPIO_PAD_fm[184];

// ----- Blif Benchmark output odata_4_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[375] -----
	assign odata_4_33_[0] = gfpga_pad_GPIO_PAD_fm[375];

// ----- Blif Benchmark output odata_4_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[444] -----
	assign odata_4_34_[0] = gfpga_pad_GPIO_PAD_fm[444];

// ----- Blif Benchmark output ovalid_4 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[22] -----
	assign ovalid_4[0] = gfpga_pad_GPIO_PAD_fm[22];

// ----- Blif Benchmark output ovch_4 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[96] -----
	assign ovch_4[0] = gfpga_pad_GPIO_PAD_fm[96];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD_fm[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[76] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[80] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[84] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[85] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[90] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[91] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[147] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[148] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[149] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[150] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[152] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[153] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[154] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[156] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[164] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[172] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[224] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[225] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[226] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[227] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[234] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[235] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[237] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[239] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[240] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[241] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[242] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[243] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[245] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[247] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[248] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[250] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[251] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[255] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[256] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[257] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[261] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[262] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[276] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[311] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[314] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[315] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[316] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[317] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[319] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[320] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[324] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[325] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[332] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[334] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[347] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[412] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[415] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
// ----- Begin assign bitstream to configuration memories -----
initial begin
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_1__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_2__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_4__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_4__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_5__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_5__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_6__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_6__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_6__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_7__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_7__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_8__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_8__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_8__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_9__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_9__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_10__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_10__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__7_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__8_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__9_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_10__10_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_8__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_9__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_10__11_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__10_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__9_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_11__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_10__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_9__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_8__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__9_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__10_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_190.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_190.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_80.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_80.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_104.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_104.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_120.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__1_.mem_top_track_120.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__1_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_102.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__1_.mem_right_track_102.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__1_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_154.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_154.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_156.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_156.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_208.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__1_.mem_right_track_208.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_145.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_145.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__2_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_66.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_66.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_112.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_112.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_146.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_146.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_154.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_154.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_156.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_156.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_186.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_186.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_200.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_200.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_209.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_209.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__3_.mem_top_track_72.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_top_track_72.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_112.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_top_track_112.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_152.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_152.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_160.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_160.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_200.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_top_track_200.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_138.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_138.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_153.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_169.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_169.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_72.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_72.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_128.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_128.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_184.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_172.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_172.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_72.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_72.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_160.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_160.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_192.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_90.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__5_.mem_right_track_90.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__5_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_180.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__5_.mem_right_track_180.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__5_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_0.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_0.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_8.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__6_.mem_top_track_8.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_48.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_48.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_64.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__6_.mem_top_track_64.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__6_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_80.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__6_.mem_top_track_80.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__6_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_152.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_152.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_192.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__6_.mem_top_track_192.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_82.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_82.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_108.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_108.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_105.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_137.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_137.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_161.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_161.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_177.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_177.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_24.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_32.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__7_.mem_top_track_32.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__7_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_128.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__7_.mem_top_track_128.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__7_.mem_top_track_136.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_0__7_.mem_top_track_136.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_0__7_.mem_top_track_144.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_144.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_176.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_176.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_200.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_84.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_84.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_92.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_92.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_148.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_148.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_154.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_154.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_200.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_200.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_25.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_41.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_41.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_49.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_49.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_137.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_209.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_209.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__8_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_16.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_32.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_32.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_40.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_40.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_36.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__8_.mem_right_track_36.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__8_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_58.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__8_.mem_right_track_58.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__8_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_98.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__8_.mem_right_track_98.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__8_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_148.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__8_.mem_right_track_148.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__8_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_160.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__8_.mem_right_track_160.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__8_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_168.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_168.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_65.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_105.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_88.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__9_.mem_top_track_88.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__9_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_54.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_54.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_176.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_176.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_186.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_186.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_202.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__9_.mem_right_track_202.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__9_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_25.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_153.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__9_.mem_bottom_track_153.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__9_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_201.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__9_.mem_bottom_track_201.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_2.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__10_.mem_right_track_2.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__10_.mem_right_track_4.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_4.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_26.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__10_.mem_right_track_26.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__10_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_62.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_62.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_84.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_84.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_150.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_150.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_172.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__10_.mem_right_track_172.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__10_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_188.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__10_.mem_right_track_188.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__10_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_right_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_right_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_141.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__10_.mem_bottom_track_141.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_136.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_top_track_136.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_164.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_top_track_164.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_120.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_right_track_120.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_152.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_152.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_80.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__1_.mem_top_track_80.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_96.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_104.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__1_.mem_top_track_104.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__1_.mem_top_track_112.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_top_track_112.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_top_track_120.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_top_track_120.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_88.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_88.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_104.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__2_.mem_top_track_104.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_176.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__2_.mem_top_track_176.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_128.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_128.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_176.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__2_.mem_right_track_176.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__2_.mem_right_track_184.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__2_.mem_right_track_184.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__2_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_161.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_left_track_161.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_136.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_136.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_105.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_105.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_105.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_left_track_105.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_129.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__3_.mem_left_track_129.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_201.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__3_.mem_left_track_201.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__3_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_128.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__4_.mem_top_track_128.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_88.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__4_.mem_right_track_88.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__4_.mem_right_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_89.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_89.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_177.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_177.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_80.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__5_.mem_right_track_80.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__5_.mem_right_track_88.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__5_.mem_right_track_88.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_168.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__6_.mem_top_track_168.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_97.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_97.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_113.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__6_.mem_left_track_113.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_185.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__6_.mem_left_track_185.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_17.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_40.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__8_.mem_top_track_40.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_120.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__8_.mem_right_track_120.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_25.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__8_.mem_left_track_25.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_48.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_48.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_80.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__9_.mem_right_track_80.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_112.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_160.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__9_.mem_right_track_160.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_65.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__9_.mem_bottom_track_65.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__9_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__9_.mem_bottom_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_72.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_184.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_13.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__10_.mem_bottom_track_13.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_35.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__10_.mem_bottom_track_35.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_159.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__10_.mem_bottom_track_159.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_145.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__10_.mem_left_track_145.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__10_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_66.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_top_track_66.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_top_track_68.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_68.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_96.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_top_track_96.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_144.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_top_track_144.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_160.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_160.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_89.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_185.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_left_track_185.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_88.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_top_track_88.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_120.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__1_.mem_top_track_120.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_168.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_right_track_168.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_184.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_184.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_193.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_193.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_left_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_left_track_121.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_193.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_left_track_193.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_80.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_top_track_80.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_104.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_top_track_104.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_128.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_top_track_128.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_top_track_136.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_top_track_136.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_top_track_144.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_top_track_144.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_160.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_top_track_160.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_184.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_top_track_184.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_200.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_top_track_200.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__2_.mem_right_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_120.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_120.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_136.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_right_track_136.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_right_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_168.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_168.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_192.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_192.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_208.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_right_track_208.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_73.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_73.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_129.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_129.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_120.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_right_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_144.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__3_.mem_right_track_144.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_168.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__3_.mem_right_track_168.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_192.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_192.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_113.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_113.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__3_.mem_left_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_177.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__3_.mem_left_track_177.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_96.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__4_.mem_top_track_96.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_184.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__4_.mem_top_track_184.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_88.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__4_.mem_right_track_88.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_144.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_right_track_144.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_176.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__4_.mem_right_track_176.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_200.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__4_.mem_right_track_200.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_153.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_153.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_81.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_96.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__5_.mem_top_track_96.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_168.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_top_track_168.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_80.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_right_track_80.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_120.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__5_.mem_right_track_120.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_136.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_right_track_136.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_right_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_right_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_right_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_184.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__5_.mem_right_track_184.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_80.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__6_.mem_top_track_80.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__6_.mem_right_track_72.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__6_.mem_right_track_72.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__6_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_96.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__6_.mem_right_track_96.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__6_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_120.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__6_.mem_right_track_120.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__6_.mem_right_track_128.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__6_.mem_right_track_128.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_144.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_right_track_144.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_right_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__6_.mem_right_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__6_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_192.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_right_track_192.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_right_track_200.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__6_.mem_right_track_200.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_81.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_81.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_97.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_97.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_121.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_121.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_161.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_161.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_169.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_169.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_177.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_177.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_185.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_8.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__7_.mem_top_track_8.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_32.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__7_.mem_top_track_32.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_128.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__7_.mem_top_track_128.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__7_.mem_top_track_136.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__7_.mem_top_track_136.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_8.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__7_.mem_right_track_8.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_24.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__7_.mem_right_track_24.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_104.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__7_.mem_right_track_104.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_41.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_41.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_137.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_137.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_9.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_33.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__7_.mem_left_track_33.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__7_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_89.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__7_.mem_left_track_89.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_8.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__8_.mem_right_track_8.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__8_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_24.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__8_.mem_right_track_24.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__8_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_48.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__8_.mem_right_track_48.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_160.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__8_.mem_right_track_160.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__8_.mem_right_track_168.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__8_.mem_right_track_168.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_25.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_25.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_73.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_73.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_81.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_81.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_137.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_137.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_177.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_177.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__8_.mem_left_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_16.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__9_.mem_top_track_16.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_104.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__9_.mem_top_track_104.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_152.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__9_.mem_top_track_152.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_184.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_0.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__9_.mem_right_track_0.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_128.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__9_.mem_right_track_128.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_160.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__9_.mem_right_track_160.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__9_.mem_bottom_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__9_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_129.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__9_.mem_bottom_track_129.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__9_.mem_bottom_track_137.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__9_.mem_bottom_track_137.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__9_.mem_left_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_185.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__9_.mem_left_track_185.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__9_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__10_.mem_right_track_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_32.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_88.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_128.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_152.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_3.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_3.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_19.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_19.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_41.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_41.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_45.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_45.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_bottom_track_209.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__10_.mem_bottom_track_209.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_73.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_73.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_97.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__10_.mem_left_track_97.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_153.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_185.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__10_.mem_left_track_185.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__10_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_18.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_top_track_18.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_116.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_top_track_116.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_88.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_104.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_104.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_144.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_right_track_144.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_73.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_left_track_73.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_177.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_left_track_177.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__1_.mem_top_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__1_.mem_top_track_80.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_80.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_120.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__1_.mem_top_track_120.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_152.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__1_.mem_top_track_152.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_152.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__1_.mem_right_track_152.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_168.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__1_.mem_right_track_168.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_200.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_right_track_200.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_201.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_left_track_201.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_80.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__2_.mem_top_track_80.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__2_.mem_top_track_88.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_top_track_88.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_112.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_top_track_112.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_144.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__2_.mem_top_track_144.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__2_.mem_top_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__2_.mem_top_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_192.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_3__2_.mem_top_track_192.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_3__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_136.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__2_.mem_right_track_136.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_192.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__2_.mem_right_track_192.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__2_.mem_right_track_200.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__2_.mem_right_track_200.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__2_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_169.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_169.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_121.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__2_.mem_left_track_121.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_201.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__2_.mem_left_track_201.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_200.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__3_.mem_top_track_200.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_104.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_right_track_104.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_144.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__3_.mem_right_track_144.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__3_.mem_right_track_152.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_right_track_152.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_201.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_201.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_81.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__3_.mem_left_track_81.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_160.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_top_track_160.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_128.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__4_.mem_right_track_128.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_144.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__4_.mem_right_track_144.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_right_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_right_track_168.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_right_track_168.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_209.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_209.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_161.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__4_.mem_left_track_161.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__5_.mem_top_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__5_.mem_top_track_80.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__5_.mem_top_track_80.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_128.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__5_.mem_top_track_128.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_152.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__5_.mem_top_track_152.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_184.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__5_.mem_top_track_184.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_200.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__5_.mem_top_track_200.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_80.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__5_.mem_right_track_80.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_96.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__5_.mem_right_track_96.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_128.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__5_.mem_right_track_128.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_144.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__5_.mem_right_track_144.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__5_.mem_right_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__5_.mem_right_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__5_.mem_right_track_160.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__5_.mem_right_track_160.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_184.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__5_.mem_right_track_184.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__5_.mem_right_track_192.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__5_.mem_right_track_192.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__5_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_104.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__6_.mem_top_track_104.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__6_.mem_right_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__6_.mem_right_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__6_.mem_right_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__6_.mem_right_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__6_.mem_right_track_88.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__6_.mem_right_track_88.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__6_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_128.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_128.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__6_.mem_right_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__6_.mem_right_track_152.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__6_.mem_right_track_152.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__6_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_176.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__6_.mem_right_track_176.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_192.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__6_.mem_right_track_192.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__6_.mem_right_track_200.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_73.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_73.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_89.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_89.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_113.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_113.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_137.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_161.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_169.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_185.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_177.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__6_.mem_left_track_177.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__6_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_120.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__7_.mem_top_track_120.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_144.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__7_.mem_right_track_144.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_41.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_41.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_65.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_65.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_145.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_145.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_41.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__7_.mem_left_track_41.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_89.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__7_.mem_left_track_89.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_8.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__8_.mem_top_track_8.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__8_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_152.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__8_.mem_right_track_152.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__8_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_65.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__8_.mem_bottom_track_65.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_56.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__9_.mem_top_track_56.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__9_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_184.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__9_.mem_top_track_184.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_64.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__9_.mem_right_track_64.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_80.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__9_.mem_right_track_80.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_144.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__9_.mem_right_track_144.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__9_.mem_right_track_152.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__9_.mem_right_track_152.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__9_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_161.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__9_.mem_bottom_track_161.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_193.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_3__9_.mem_bottom_track_193.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_3__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_41.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__9_.mem_left_track_41.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_65.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__9_.mem_left_track_65.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_81.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__9_.mem_left_track_81.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_112.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_128.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_144.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_192.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__10_.mem_right_track_192.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_139.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__10_.mem_bottom_track_139.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__10_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__10_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_49.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_49.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_73.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__10_.mem_left_track_73.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__10_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_97.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__10_.mem_left_track_97.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_113.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__10_.mem_left_track_113.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_145.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__10_.mem_left_track_145.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__10_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_136.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__0_.mem_right_track_136.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_184.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__0_.mem_right_track_184.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_89.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__0_.mem_left_track_89.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_129.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_145.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__0_.mem_left_track_145.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_185.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__0_.mem_left_track_185.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__0_.mem_left_track_193.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__0_.mem_left_track_193.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_80.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_top_track_80.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_96.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_112.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_136.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_top_track_136.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_top_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_top_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_top_track_152.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_top_track_152.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_192.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_top_track_192.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_32.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_right_track_32.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_56.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_right_track_56.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__1_.mem_right_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_128.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_right_track_128.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_left_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_104.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__2_.mem_top_track_104.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_152.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__2_.mem_top_track_152.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_8.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__2_.mem_right_track_8.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_40.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__2_.mem_right_track_40.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_56.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__2_.mem_right_track_56.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_80.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__2_.mem_right_track_80.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_176.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__2_.mem_right_track_176.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__2_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_169.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_169.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_113.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_113.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_201.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__2_.mem_left_track_201.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_80.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__3_.mem_top_track_80.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__3_.mem_top_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_160.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_96.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_104.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__3_.mem_right_track_104.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_120.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__3_.mem_right_track_120.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_168.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__3_.mem_right_track_168.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_184.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__3_.mem_right_track_184.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_177.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_177.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__3_.mem_left_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_209.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_left_track_209.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_152.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__4_.mem_top_track_152.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_112.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__4_.mem_right_track_112.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_184.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__4_.mem_right_track_184.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_105.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_105.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_161.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_161.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_185.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_185.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__5_.mem_top_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_200.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__5_.mem_top_track_200.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__5_.mem_right_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_24.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__5_.mem_right_track_24.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__5_.mem_right_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_88.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__5_.mem_right_track_88.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_120.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__5_.mem_right_track_120.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__5_.mem_right_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_160.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__5_.mem_right_track_160.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_right_track_200.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__5_.mem_right_track_200.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__5_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_121.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_121.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_145.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_145.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_193.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_193.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__6_.mem_top_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_0.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__6_.mem_right_track_0.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_24.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_32.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__6_.mem_right_track_32.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__6_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_48.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__6_.mem_right_track_48.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__6_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_64.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__6_.mem_right_track_64.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__6_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__6_.mem_right_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__6_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__6_.mem_right_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__6_.mem_right_track_168.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__6_.mem_right_track_168.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__6_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_right_track_200.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__6_.mem_right_track_200.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_73.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_73.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_105.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_105.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_177.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_177.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_193.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_193.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_153.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__6_.mem_left_track_153.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_73.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_73.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_193.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_193.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_209.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_209.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_4__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_0.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__8_.mem_top_track_0.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__8_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_0.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__8_.mem_right_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_88.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__8_.mem_right_track_88.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__8_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_153.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__8_.mem_bottom_track_153.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__8_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_128.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__9_.mem_right_track_128.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_176.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__9_.mem_right_track_176.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__9_.mem_bottom_track_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_17.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__9_.mem_bottom_track_17.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_169.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__9_.mem_bottom_track_169.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_128.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_57.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_57.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_67.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_67.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_83.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_83.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_97.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_97.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_9.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__10_.mem_left_track_9.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__10_.mem_left_track_17.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_17.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_25.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__10_.mem_left_track_25.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_105.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__10_.mem_left_track_105.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__10_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_193.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__10_.mem_left_track_193.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_50.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_5__0_.mem_top_track_50.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_5__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_64.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_5__0_.mem_top_track_64.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_5__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_100.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__0_.mem_top_track_100.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_108.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__0_.mem_top_track_108.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_180.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__0_.mem_top_track_180.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_72.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_5__0_.mem_right_track_72.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_5__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_96.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__0_.mem_right_track_96.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_120.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_right_track_208.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_5__0_.mem_right_track_208.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_5__0_.mem_left_track_1.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__0_.mem_left_track_1.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_81.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_89.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__0_.mem_left_track_89.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_169.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__0_.mem_left_track_169.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_16.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__1_.mem_top_track_16.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_136.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_200.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_136.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__1_.mem_right_track_136.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_121.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_121.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_41.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__1_.mem_left_track_41.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_89.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__1_.mem_left_track_89.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__1_.mem_left_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_8.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__2_.mem_top_track_8.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_24.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__2_.mem_top_track_24.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__2_.mem_top_track_32.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_56.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__2_.mem_top_track_56.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__2_.mem_top_track_64.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__2_.mem_top_track_64.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_96.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__2_.mem_top_track_96.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_176.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__2_.mem_top_track_176.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_192.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_5__2_.mem_top_track_192.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_5__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_24.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__2_.mem_right_track_24.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__2_.mem_right_track_32.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__2_.mem_right_track_32.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_56.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__2_.mem_right_track_56.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_72.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__2_.mem_right_track_72.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_88.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__2_.mem_right_track_88.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__2_.mem_right_track_96.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__2_.mem_right_track_96.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__2_.mem_right_track_104.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__2_.mem_right_track_104.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_120.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__2_.mem_right_track_120.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_152.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__2_.mem_right_track_152.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_81.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_81.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_161.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_161.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_177.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_177.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_33.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__2_.mem_left_track_33.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_81.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__2_.mem_left_track_81.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_113.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__2_.mem_left_track_113.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_185.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__2_.mem_left_track_185.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__2_.mem_left_track_201.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__2_.mem_left_track_201.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_24.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_5__3_.mem_top_track_24.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_5__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_56.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__3_.mem_top_track_56.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__3_.mem_top_track_64.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__3_.mem_top_track_64.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_96.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__3_.mem_top_track_96.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__3_.mem_top_track_104.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__3_.mem_top_track_104.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__3_.mem_top_track_112.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__3_.mem_top_track_112.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_128.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_136.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_144.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__3_.mem_top_track_144.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_176.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__3_.mem_top_track_176.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__3_.mem_right_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__3_.mem_right_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_112.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_144.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_168.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__3_.mem_right_track_168.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_right_track_208.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_5__3_.mem_right_track_208.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_25.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_25.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_81.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_81.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__3_.mem_left_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_33.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__3_.mem_left_track_33.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_57.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__3_.mem_left_track_57.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_153.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__3_.mem_left_track_153.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_201.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__3_.mem_left_track_201.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_8.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__4_.mem_top_track_8.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_32.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__4_.mem_top_track_32.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__4_.mem_top_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__4_.mem_top_track_64.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_72.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__4_.mem_top_track_72.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__4_.mem_top_track_80.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__4_.mem_top_track_80.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_96.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__4_.mem_top_track_96.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_136.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__4_.mem_top_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_176.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__4_.mem_top_track_176.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__4_.mem_top_track_184.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__4_.mem_top_track_184.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_top_track_200.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_5__4_.mem_top_track_200.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_5__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_40.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_64.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__4_.mem_right_track_64.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_136.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__4_.mem_right_track_136.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_160.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__4_.mem_right_track_160.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_184.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_right_track_208.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_5__4_.mem_right_track_208.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_209.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_209.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__4_.mem_left_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_41.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__4_.mem_left_track_41.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_113.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__4_.mem_left_track_113.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_137.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__4_.mem_left_track_137.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_177.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__4_.mem_left_track_177.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_top_track_0.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_top_track_0.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_top_track_8.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_16.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_top_track_16.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_top_track_24.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_top_track_24.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_top_track_32.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_top_track_32.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_top_track_40.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_top_track_40.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_top_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_top_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_top_track_56.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_top_track_56.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_top_track_64.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_top_track_64.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_top_track_72.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_top_track_72.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_top_track_80.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_top_track_80.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_top_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_96.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__5_.mem_top_track_96.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__5_.mem_top_track_104.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_top_track_104.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_top_track_112.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__5_.mem_top_track_112.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__5_.mem_top_track_120.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_top_track_120.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_top_track_128.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_136.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__5_.mem_top_track_136.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__5_.mem_top_track_144.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_top_track_144.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_top_track_152.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__5_.mem_top_track_152.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__5_.mem_top_track_160.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_top_track_160.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_top_track_168.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_top_track_168.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_top_track_176.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__5_.mem_top_track_176.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__5_.mem_top_track_184.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_top_track_184.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_top_track_192.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__5_.mem_top_track_192.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__5_.mem_top_track_200.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_top_track_200.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_top_track_208.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_top_track_208.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_right_track_0.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_right_track_0.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_right_track_8.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_8.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_24.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_right_track_24.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_32.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_32.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_40.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_40.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_right_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_right_track_56.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_56.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_64.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_right_track_64.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_72.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_72.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_right_track_80.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_right_track_80.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_right_track_88.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_right_track_88.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_right_track_96.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_96.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_104.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_104.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_right_track_112.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_right_track_112.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_right_track_120.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_120.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_128.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_right_track_128.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_right_track_136.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_right_track_136.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_right_track_144.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_right_track_144.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_160.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_right_track_160.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_168.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_168.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_right_track_176.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_176.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_184.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_right_track_184.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_right_track_192.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__5_.mem_right_track_192.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__5_.mem_right_track_200.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__5_.mem_right_track_200.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__5_.mem_right_track_208.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__5_.mem_right_track_208.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_33.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_33.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_81.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_81.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_201.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_201.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_209.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_209.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__5_.mem_left_track_1.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_left_track_1.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_left_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__5_.mem_left_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_97.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__5_.mem_left_track_97.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__5_.mem_left_track_209.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_5__5_.mem_left_track_209.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_5__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_top_track_200.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__6_.mem_top_track_200.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_right_track_0.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_right_track_0.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_right_track_8.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_right_track_8.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_right_track_16.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_right_track_16.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_right_track_24.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_right_track_24.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_right_track_32.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_right_track_32.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_right_track_40.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_40.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_48.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_right_track_48.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_right_track_56.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_56.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_64.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_right_track_64.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_right_track_72.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_72.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_80.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_80.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_88.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_right_track_88.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_right_track_96.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_right_track_96.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_right_track_104.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_104.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_112.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_112.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_120.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_right_track_120.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_right_track_128.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_right_track_128.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_right_track_136.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_right_track_136.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_right_track_144.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_right_track_144.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_right_track_152.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_right_track_152.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_right_track_160.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_right_track_160.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_right_track_168.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_right_track_168.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_right_track_176.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_176.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_184.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_right_track_184.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_right_track_192.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_right_track_192.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_right_track_200.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__6_.mem_right_track_200.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__6_.mem_right_track_208.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_right_track_208.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_9.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_9.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_17.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_17.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_25.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_25.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_33.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_33.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_41.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_41.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_49.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_49.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_57.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_57.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_65.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_65.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_73.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_73.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_81.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_81.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_89.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_89.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_105.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_105.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_113.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_113.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_121.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_121.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_129.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_129.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_137.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_137.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_145.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_145.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_153.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_153.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_161.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_161.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_169.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_169.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_177.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_177.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_185.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_185.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_193.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_193.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_201.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_201.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_209.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_209.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__6_.mem_left_track_1.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_left_track_1.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_left_track_9.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_left_track_9.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_57.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__6_.mem_left_track_57.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__6_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__6_.mem_left_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__6_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_105.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__6_.mem_left_track_105.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_177.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__6_.mem_left_track_177.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__6_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_0.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__7_.mem_right_track_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_72.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__7_.mem_right_track_72.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_168.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__7_.mem_right_track_168.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_192.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__7_.mem_right_track_192.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_41.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_41.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_81.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_81.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_121.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_121.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_65.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__7_.mem_left_track_65.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__7_.mem_left_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_40.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__8_.mem_right_track_40.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__8_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_88.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__8_.mem_right_track_88.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__8_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_112.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__8_.mem_right_track_112.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__8_.mem_right_track_120.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__8_.mem_right_track_120.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_160.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__8_.mem_right_track_160.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_184.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__8_.mem_right_track_184.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__8_.mem_right_track_192.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__8_.mem_right_track_192.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_25.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_25.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_41.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_41.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_57.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_81.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_81.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_113.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_113.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_137.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_137.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_153.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_153.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_161.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_161.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_49.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__8_.mem_left_track_49.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_64.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__9_.mem_top_track_64.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_120.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__9_.mem_top_track_120.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_152.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__9_.mem_top_track_152.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__9_.mem_right_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__9_.mem_right_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__9_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_120.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__9_.mem_right_track_120.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__9_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_136.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__9_.mem_right_track_136.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__9_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__9_.mem_right_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__9_.mem_right_track_160.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__9_.mem_right_track_160.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_184.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__9_.mem_right_track_184.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_57.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_57.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_73.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_73.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_153.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_153.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_161.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_161.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_177.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_177.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_185.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_185.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_193.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_193.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_5__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_65.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_5__9_.mem_left_track_65.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_5__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_137.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__9_.mem_left_track_137.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_177.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__9_.mem_left_track_177.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__9_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_193.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_5__9_.mem_left_track_193.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_5__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_24.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_5__10_.mem_right_track_24.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_5__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_48.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_72.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_88.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_109.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_5__10_.mem_bottom_track_109.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_5__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_117.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_5__10_.mem_bottom_track_117.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_5__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_189.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_5__10_.mem_bottom_track_189.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_5__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_49.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_5__10_.mem_left_track_49.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_5__10_.mem_left_track_57.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_5__10_.mem_left_track_57.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_5__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_73.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__10_.mem_left_track_73.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__10_.mem_left_track_81.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__10_.mem_left_track_81.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_169.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__10_.mem_left_track_169.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_185.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_5__10_.mem_left_track_185.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_5__10_.mem_left_track_193.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_5__10_.mem_left_track_193.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_5__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_5__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_92.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_96.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_108.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_6__0_.mem_top_track_108.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_6__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_118.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_6__0_.mem_top_track_118.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_6__0_.mem_top_track_120.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_148.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_152.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_170.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_6__0_.mem_top_track_170.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_6__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_168.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__0_.mem_right_track_168.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_1.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_6__0_.mem_left_track_1.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_6__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_17.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_73.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__0_.mem_left_track_73.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_89.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__0_.mem_left_track_89.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_153.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__0_.mem_left_track_153.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_169.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_left_track_201.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_6__0_.mem_left_track_201.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_6__0_.mem_left_track_209.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__0_.mem_left_track_209.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_32.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__1_.mem_top_track_32.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_72.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__1_.mem_top_track_72.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__1_.mem_top_track_80.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_80.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_top_track_208.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__1_.mem_top_track_208.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_24.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__1_.mem_right_track_24.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_72.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__1_.mem_right_track_72.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__1_.mem_right_track_80.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__1_.mem_right_track_80.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_right_track_208.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_6__1_.mem_right_track_208.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_169.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_169.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_33.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__1_.mem_left_track_33.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_57.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__1_.mem_left_track_57.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_121.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__1_.mem_left_track_121.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_8.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__2_.mem_top_track_8.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__2_.mem_top_track_16.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_6__2_.mem_top_track_16.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_6__2_.mem_top_track_24.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_6__2_.mem_top_track_24.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_6__2_.mem_top_track_32.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_56.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_96.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__2_.mem_top_track_96.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_112.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_top_track_112.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_144.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__2_.mem_top_track_144.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_112.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__2_.mem_right_track_112.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__2_.mem_right_track_120.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_right_track_120.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_136.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_right_track_136.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_160.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_right_track_160.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_176.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_right_track_176.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_right_track_184.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_right_track_184.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_right_track_192.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_right_track_192.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_17.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_17.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_25.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_25.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_49.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_49.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_57.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_57.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_161.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_161.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_209.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_209.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__2_.mem_left_track_1.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__2_.mem_left_track_1.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__2_.mem_left_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__2_.mem_left_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__2_.mem_left_track_17.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__2_.mem_left_track_17.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__2_.mem_left_track_25.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__2_.mem_left_track_25.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_57.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_left_track_57.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_73.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_left_track_73.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_left_track_81.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_left_track_81.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__2_.mem_left_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__2_.mem_left_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__2_.mem_left_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_169.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__2_.mem_left_track_169.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_185.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__2_.mem_left_track_185.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__3_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_24.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_6__3_.mem_top_track_24.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_6__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_56.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__3_.mem_top_track_56.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_72.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__3_.mem_top_track_72.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__3_.mem_top_track_80.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__3_.mem_top_track_80.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_96.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__3_.mem_top_track_96.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__3_.mem_top_track_104.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__3_.mem_top_track_104.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__3_.mem_top_track_112.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__3_.mem_top_track_112.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__3_.mem_top_track_120.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__3_.mem_top_track_120.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_136.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__3_.mem_top_track_136.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_168.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__3_.mem_top_track_168.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__3_.mem_top_track_176.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__3_.mem_top_track_176.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_48.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_120.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__3_.mem_right_track_120.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_9.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_9.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_65.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_65.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_145.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_145.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_209.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_209.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_6__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_49.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__3_.mem_left_track_49.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_89.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__3_.mem_left_track_89.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__3_.mem_left_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_129.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_161.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__3_.mem_left_track_161.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__3_.mem_left_track_169.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__3_.mem_left_track_169.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__3_.mem_left_track_177.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__3_.mem_left_track_177.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_201.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__3_.mem_left_track_201.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_0.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__4_.mem_top_track_0.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__4_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__4_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_24.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__4_.mem_top_track_24.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__4_.mem_top_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_56.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__4_.mem_top_track_56.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_88.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__4_.mem_top_track_88.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_128.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__4_.mem_top_track_128.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_160.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__4_.mem_top_track_160.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__4_.mem_top_track_168.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_184.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_192.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_6__4_.mem_top_track_192.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_6__4_.mem_top_track_200.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_6__4_.mem_top_track_200.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_6__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_64.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_136.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_9.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__4_.mem_left_track_9.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__4_.mem_left_track_17.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_25.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__4_.mem_left_track_25.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_41.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_49.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__4_.mem_left_track_49.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_65.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__4_.mem_left_track_65.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_105.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__4_.mem_left_track_105.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_137.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__4_.mem_left_track_137.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__4_.mem_left_track_209.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_6__4_.mem_left_track_209.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_6__5_.mem_top_track_0.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_8.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_16.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_top_track_16.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_top_track_24.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__5_.mem_top_track_24.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__5_.mem_top_track_32.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_top_track_32.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_top_track_40.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__5_.mem_top_track_40.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__5_.mem_top_track_48.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_top_track_48.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_top_track_56.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_top_track_56.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_top_track_64.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_top_track_64.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_top_track_72.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__5_.mem_top_track_72.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__5_.mem_top_track_80.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_top_track_80.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_top_track_88.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_top_track_88.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_top_track_96.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_top_track_96.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_top_track_104.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_top_track_104.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_top_track_112.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_top_track_112.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_top_track_120.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_top_track_120.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_top_track_128.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_top_track_128.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_top_track_136.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_top_track_136.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_top_track_144.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_top_track_144.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_top_track_152.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_top_track_152.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_top_track_160.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_168.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_top_track_168.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_top_track_176.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_top_track_176.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_top_track_184.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_top_track_184.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_192.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_top_track_192.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_top_track_200.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__5_.mem_top_track_200.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__5_.mem_top_track_208.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_0.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_6__5_.mem_right_track_0.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_6__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_56.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_right_track_56.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_152.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_17.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_17.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_65.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_65.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_89.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_89.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_185.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_185.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_201.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_201.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__5_.mem_left_track_1.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_left_track_1.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_left_track_9.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_left_track_9.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_left_track_17.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_17.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_25.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__5_.mem_left_track_25.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__5_.mem_left_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_41.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_left_track_41.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_left_track_49.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_left_track_49.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_left_track_57.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_57.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_65.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__5_.mem_left_track_65.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__5_.mem_left_track_73.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__5_.mem_left_track_73.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__5_.mem_left_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_89.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_left_track_89.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_left_track_97.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__5_.mem_left_track_97.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__5_.mem_left_track_105.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_left_track_105.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_left_track_113.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_left_track_113.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_left_track_121.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_left_track_121.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_left_track_129.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_left_track_129.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_left_track_137.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__5_.mem_left_track_137.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__5_.mem_left_track_145.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_145.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_153.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_left_track_153.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__5_.mem_left_track_161.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_161.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_169.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_169.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_177.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__5_.mem_left_track_177.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__5_.mem_left_track_185.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__5_.mem_left_track_185.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__5_.mem_left_track_193.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__5_.mem_left_track_193.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__5_.mem_left_track_201.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__5_.mem_left_track_201.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__5_.mem_left_track_209.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__5_.mem_left_track_209.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_24.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__6_.mem_top_track_24.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_120.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_top_track_120.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_32.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_right_track_32.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_right_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_104.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_right_track_104.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_152.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_right_track_152.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__6_.mem_right_track_208.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__6_.mem_right_track_208.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_9.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_9.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_17.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_17.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_25.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_25.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_41.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_41.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_49.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_49.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_57.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_57.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_65.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_65.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_73.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_73.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_81.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_81.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_89.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_89.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_105.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_105.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_121.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_121.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_129.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_129.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_137.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_137.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_145.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_145.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_161.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_161.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_169.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_169.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_177.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_177.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_185.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_185.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_193.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_193.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_201.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_201.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_209.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_209.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_1.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_left_track_1.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_left_track_9.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_9.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_left_track_17.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_17.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_left_track_25.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_25.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_left_track_33.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_left_track_33.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_left_track_41.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_left_track_41.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_left_track_49.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_left_track_49.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_left_track_57.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_57.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_left_track_65.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_left_track_65.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_left_track_73.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_left_track_73.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_left_track_81.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_left_track_81.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_left_track_89.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_89.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_left_track_97.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_left_track_97.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_left_track_105.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_left_track_105.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_left_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_left_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_left_track_121.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_left_track_121.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_left_track_129.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_left_track_129.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_left_track_137.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__6_.mem_left_track_137.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__6_.mem_left_track_145.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_left_track_145.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_left_track_153.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__6_.mem_left_track_153.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__6_.mem_left_track_161.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__6_.mem_left_track_161.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__6_.mem_left_track_169.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_169.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_left_track_177.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_left_track_177.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_left_track_185.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_left_track_185.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_left_track_193.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__6_.mem_left_track_193.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__6_.mem_left_track_201.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__6_.mem_left_track_201.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__6_.mem_left_track_209.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__6_.mem_left_track_209.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_96.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__7_.mem_right_track_96.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__7_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_120.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__7_.mem_right_track_120.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_192.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__7_.mem_right_track_192.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_1.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_1.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_41.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_41.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_97.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_97.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_137.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_137.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_17.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_6__7_.mem_left_track_17.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_6__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_41.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__7_.mem_left_track_41.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__7_.mem_left_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__7_.mem_left_track_121.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__7_.mem_left_track_121.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_137.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__7_.mem_left_track_137.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_161.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__7_.mem_left_track_161.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_185.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__7_.mem_left_track_185.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__8_.mem_top_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__8_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_40.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__8_.mem_right_track_40.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__8_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_64.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__8_.mem_right_track_64.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_112.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__8_.mem_right_track_112.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__8_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_57.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_57.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_137.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_137.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_145.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_145.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_153.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_153.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_169.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_169.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_1.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__8_.mem_left_track_1.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__8_.mem_left_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__8_.mem_left_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_49.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__8_.mem_left_track_49.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_145.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__8_.mem_left_track_145.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_6__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_48.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__9_.mem_right_track_48.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_104.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__9_.mem_right_track_104.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_128.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__9_.mem_right_track_128.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_160.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_6__9_.mem_right_track_160.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_6__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_1.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_1.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_9.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_9.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_25.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_25.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_33.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_33.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_41.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_41.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_73.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_73.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_121.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_121.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_137.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_137.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_185.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_185.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_bottom_track_201.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_201.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_209.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_6__9_.mem_bottom_track_209.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_6__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_25.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_6__9_.mem_left_track_25.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_6__9_.mem_left_track_33.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_6__9_.mem_left_track_33.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_6__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_81.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__9_.mem_left_track_81.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_6__9_.mem_left_track_89.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__9_.mem_left_track_89.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__9_.mem_left_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_6__9_.mem_left_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_6__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_56.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_80.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_6__10_.mem_right_track_80.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_6__10_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_184.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_99.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_6__10_.mem_bottom_track_99.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_6__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_25.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_6__10_.mem_left_track_25.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_6__10_.mem_left_track_33.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_6__10_.mem_left_track_33.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_6__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_81.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_6__10_.mem_left_track_81.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_6__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_6__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_32.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_32.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_40.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__0_.mem_top_track_40.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_72.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__0_.mem_top_track_72.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_80.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__0_.mem_top_track_80.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__0_.mem_top_track_82.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__0_.mem_top_track_82.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_146.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__0_.mem_top_track_146.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_24.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__0_.mem_right_track_24.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_40.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__0_.mem_right_track_40.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_64.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__0_.mem_right_track_64.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_88.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__0_.mem_right_track_88.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__0_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_49.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_65.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_7__0_.mem_left_track_65.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_7__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_81.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__0_.mem_left_track_81.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_113.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_161.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__0_.mem_left_track_161.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_160.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_168.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__1_.mem_top_track_168.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_192.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__1_.mem_top_track_192.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_56.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__1_.mem_right_track_56.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_105.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_105.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_201.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_201.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_1.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__1_.mem_left_track_1.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_81.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__1_.mem_left_track_81.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_97.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__1_.mem_left_track_97.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_121.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__1_.mem_left_track_121.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_16.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_7__2_.mem_top_track_16.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_7__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_112.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__2_.mem_top_track_112.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__2_.mem_top_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_0.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_7__2_.mem_right_track_0.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_7__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_96.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_right_track_208.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_7__2_.mem_right_track_208.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_25.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_25.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_41.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_41.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_97.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_97.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_49.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__2_.mem_left_track_49.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_81.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__2_.mem_left_track_81.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_121.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__2_.mem_left_track_121.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_137.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__2_.mem_left_track_137.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_7__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_153.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__2_.mem_left_track_153.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_193.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__2_.mem_left_track_193.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_184.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__3_.mem_right_track_184.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_1.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_1.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_97.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_97.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_209.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_209.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_7__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_49.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__3_.mem_left_track_49.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__3_.mem_left_track_57.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_121.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__3_.mem_left_track_121.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__3_.mem_left_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_201.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_7__3_.mem_left_track_201.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_7__3_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_24.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_7__4_.mem_top_track_24.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_7__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__4_.mem_top_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_16.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__4_.mem_right_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_9.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_9.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_121.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_121.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_65.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__4_.mem_left_track_65.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_152.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__5_.mem_top_track_152.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_144.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__5_.mem_right_track_144.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_176.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__5_.mem_right_track_176.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_7__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_1.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_1.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_25.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_25.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_49.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_49.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_121.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_121.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_129.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_145.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__5_.mem_left_track_145.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_169.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__5_.mem_left_track_169.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__5_.mem_left_track_177.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__5_.mem_left_track_177.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_88.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__6_.mem_top_track_88.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_1.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_1.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_25.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_25.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_49.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_49.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_73.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_73.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_97.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_97.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_201.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_201.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__6_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_33.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__6_.mem_left_track_33.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__6_.mem_left_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_7__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_153.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__6_.mem_left_track_153.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_72.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_7__7_.mem_top_track_72.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_112.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__7_.mem_right_track_112.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_24.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_7__8_.mem_top_track_24.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_7__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_88.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__8_.mem_top_track_88.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_7__8_.mem_top_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_56.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__8_.mem_right_track_56.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_7__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_25.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__8_.mem_bottom_track_25.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_7__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__8_.mem_bottom_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_137.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__8_.mem_bottom_track_137.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_7__8_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_32.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__9_.mem_top_track_32.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_88.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__9_.mem_top_track_88.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_7__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_184.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_7__9_.mem_top_track_184.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_7__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_161.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__9_.mem_bottom_track_161.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__9_.mem_left_track_209.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_7__9_.mem_left_track_209.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_7__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_72.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__10_.mem_right_track_72.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_96.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_112.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_7__10_.mem_right_track_112.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_7__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_128.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_152.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_184.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_right_track_200.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__10_.mem_right_track_200.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_97.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_7__10_.mem_left_track_97.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_7__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_113.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_121.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_7__10_.mem_left_track_121.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_7__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_145.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__10_.mem_left_track_145.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__10_.mem_left_track_153.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__10_.mem_left_track_153.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_169.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__10_.mem_left_track_169.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_7__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_7__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_82.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_top_track_82.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_144.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_top_track_144.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_162.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__0_.mem_top_track_162.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_8__0_.mem_top_track_164.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_top_track_164.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_180.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__0_.mem_top_track_180.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_8__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_192.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__0_.mem_top_track_192.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_8__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_32.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_right_track_32.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_88.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_right_track_88.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_104.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_right_track_104.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_160.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_right_track_160.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_9.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_left_track_9.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_25.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_41.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__0_.mem_left_track_41.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_8__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_89.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__0_.mem_left_track_89.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_8__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_129.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_left_track_129.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_145.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__0_.mem_left_track_145.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_0.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__1_.mem_top_track_0.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__1_.mem_top_track_8.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__1_.mem_top_track_8.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_24.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__1_.mem_top_track_24.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_80.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_top_track_80.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_top_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_120.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__1_.mem_top_track_120.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_160.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__1_.mem_top_track_160.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__1_.mem_top_track_168.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_top_track_168.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_top_track_176.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_184.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_top_track_184.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_40.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_right_track_40.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_64.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_right_track_64.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__1_.mem_right_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_136.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_right_track_136.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_right_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_right_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_49.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__1_.mem_bottom_track_49.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_161.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__1_.mem_bottom_track_161.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_145.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__1_.mem_left_track_145.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_169.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__1_.mem_left_track_169.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_209.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__1_.mem_left_track_209.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__2_.mem_top_track_0.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_top_track_0.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__2_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__2_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_32.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__2_.mem_top_track_32.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_64.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__2_.mem_top_track_64.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_80.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__2_.mem_top_track_80.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_24.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__2_.mem_right_track_24.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__2_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_48.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_right_track_48.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_120.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__2_.mem_right_track_120.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_184.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_184.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_97.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_97.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_129.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_129.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_145.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_145.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_161.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_161.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_193.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_193.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_9.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__2_.mem_left_track_9.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_41.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_left_track_41.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_65.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_left_track_65.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_121.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__2_.mem_left_track_121.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_153.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__2_.mem_left_track_153.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_40.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__3_.mem_right_track_40.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_120.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_81.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_81.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_89.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_89.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_105.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_105.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_129.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_129.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_25.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_8__3_.mem_left_track_25.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_8__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_41.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__3_.mem_left_track_41.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_89.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__3_.mem_left_track_89.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_105.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__3_.mem_left_track_105.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__3_.mem_left_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__3_.mem_left_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__3_.mem_left_track_209.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__3_.mem_left_track_209.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_8__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_80.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__4_.mem_top_track_80.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__4_.mem_top_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_104.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__4_.mem_top_track_104.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_144.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__4_.mem_top_track_144.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_136.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__4_.mem_right_track_136.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_168.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__4_.mem_right_track_168.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_57.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_57.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_153.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_153.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_193.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_193.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_201.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_201.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_57.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__4_.mem_left_track_57.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_73.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__4_.mem_left_track_73.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_97.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__4_.mem_left_track_97.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_137.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_145.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__4_.mem_left_track_145.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_185.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__4_.mem_left_track_185.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__4_.mem_left_track_201.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_8__4_.mem_left_track_201.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_8__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_56.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__5_.mem_top_track_56.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_128.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__5_.mem_top_track_128.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_152.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__5_.mem_top_track_152.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__5_.mem_top_track_160.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_176.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__5_.mem_right_track_176.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_9.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_9.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_81.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_81.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_177.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_177.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_25.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__5_.mem_left_track_25.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_8__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_81.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__5_.mem_left_track_81.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_97.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__5_.mem_left_track_97.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__5_.mem_left_track_105.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__5_.mem_left_track_105.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_129.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__5_.mem_left_track_129.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_145.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__5_.mem_left_track_145.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_169.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__5_.mem_left_track_169.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__5_.mem_left_track_177.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__5_.mem_left_track_177.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__6_.mem_top_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_104.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__6_.mem_top_track_104.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_176.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__6_.mem_top_track_176.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_top_track_200.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_8__6_.mem_top_track_200.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_8__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_25.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_25.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_81.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_81.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_129.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_129.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_153.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_153.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_177.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_177.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__6_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_33.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__6_.mem_left_track_33.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_57.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__6_.mem_left_track_57.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__6_.mem_left_track_65.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__6_.mem_left_track_65.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__6_.mem_left_track_73.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__6_.mem_left_track_73.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__6_.mem_left_track_81.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__6_.mem_left_track_81.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__6_.mem_left_track_89.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__6_.mem_left_track_89.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_185.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__6_.mem_left_track_185.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_64.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__7_.mem_top_track_64.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__7_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_top_track_200.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__7_.mem_top_track_200.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_24.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__7_.mem_right_track_24.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__7_.mem_right_track_32.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__7_.mem_right_track_32.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_104.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__7_.mem_right_track_104.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_152.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__7_.mem_right_track_152.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_9.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__7_.mem_bottom_track_9.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_32.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__8_.mem_right_track_32.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__8_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_96.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__8_.mem_right_track_96.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_176.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__8_.mem_right_track_176.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_8__8_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_97.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_97.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_113.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_113.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_121.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_121.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_129.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_129.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_161.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_161.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_89.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__8_.mem_left_track_89.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__8_.mem_left_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_64.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__9_.mem_top_track_64.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_8__9_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_32.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__9_.mem_right_track_32.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_48.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_8__9_.mem_right_track_48.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_8__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_144.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__9_.mem_right_track_144.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_8__9_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_73.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_73.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_121.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_121.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_129.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_129.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_185.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_185.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_201.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_201.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_33.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__9_.mem_left_track_33.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_8__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_49.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_97.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__9_.mem_left_track_97.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_129.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__9_.mem_left_track_129.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_153.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__9_.mem_left_track_153.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_185.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__9_.mem_left_track_185.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_8__9_.mem_left_track_193.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_8__9_.mem_left_track_193.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_128.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_144.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__10_.mem_right_track_144.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_8__10_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_168.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_31.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_31.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_57.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_57.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_71.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_71.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_95.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_95.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_113.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_113.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_191.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_191.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_8__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_49.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__10_.mem_left_track_49.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_8__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_177.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__10_.mem_left_track_177.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_8__10_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_0.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_9__0_.mem_top_track_0.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_9__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_20.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_22.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_24.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_9__0_.mem_top_track_24.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_9__0_.mem_top_track_26.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_26.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_28.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_30.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_30.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_38.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_38.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_42.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_42.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_44.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_46.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_46.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_58.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_58.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_60.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_60.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_62.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_62.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_66.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_66.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_74.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_74.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_76.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_76.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_78.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_78.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_82.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_82.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_84.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_84.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_90.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_90.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_92.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_92.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_94.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_94.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_98.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_98.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_100.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_100.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_102.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_102.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_110.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_110.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_114.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_114.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_116.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_116.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_118.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_118.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_126.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_126.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_130.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_130.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_132.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_132.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_134.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_134.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_138.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_138.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_144.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_9__0_.mem_top_track_144.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_9__0_.mem_top_track_146.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_146.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_148.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_148.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_150.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_150.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_164.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_164.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_166.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_166.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_170.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_170.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_172.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_172.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_174.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_174.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_180.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_180.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_182.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_182.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_186.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_186.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_188.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_188.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_190.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_190.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_198.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_198.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_202.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_202.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_204.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_204.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_206.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_206.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_184.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_208.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_25.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_9__0_.mem_left_track_25.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_9__0_.mem_left_track_33.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_9__0_.mem_left_track_33.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_9__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_113.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_0.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__1_.mem_top_track_0.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_24.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__1_.mem_top_track_24.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__1_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_48.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_56.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__1_.mem_top_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__1_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_104.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__1_.mem_top_track_104.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_144.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__1_.mem_top_track_144.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_184.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_16.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__1_.mem_right_track_16.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_9__1_.mem_right_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_9__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_176.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_25.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__1_.mem_left_track_25.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_65.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__1_.mem_left_track_65.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_137.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__1_.mem_left_track_137.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_24.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_9__2_.mem_top_track_24.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_9__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_56.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_80.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__2_.mem_top_track_80.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__2_.mem_top_track_88.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__2_.mem_top_track_88.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_120.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__2_.mem_top_track_120.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_144.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__2_.mem_top_track_144.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_160.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__2_.mem_top_track_160.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_176.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__2_.mem_top_track_176.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_96.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__2_.mem_right_track_96.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_25.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_25.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_49.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_49.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_57.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_57.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_153.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_153.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__2_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_9.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__2_.mem_left_track_9.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__2_.mem_left_track_17.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__2_.mem_left_track_17.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__2_.mem_left_track_25.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__2_.mem_left_track_25.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__2_.mem_left_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_169.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__2_.mem_left_track_169.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_88.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__3_.mem_top_track_88.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_168.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__3_.mem_top_track_168.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_88.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_168.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__3_.mem_right_track_168.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_41.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__3_.mem_bottom_track_41.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_137.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__3_.mem_bottom_track_137.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_153.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__3_.mem_bottom_track_153.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_25.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_9__3_.mem_left_track_25.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_9__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_65.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__3_.mem_left_track_65.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__3_.mem_left_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__3_.mem_left_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__3_.mem_left_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_177.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__3_.mem_left_track_177.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__3_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__3_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_32.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__4_.mem_top_track_32.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__4_.mem_top_track_40.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__4_.mem_top_track_40.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__4_.mem_top_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_112.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__4_.mem_right_track_112.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_128.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_136.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__4_.mem_right_track_136.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__4_.mem_bottom_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_185.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_9__4_.mem_bottom_track_185.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_9__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__4_.mem_left_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__4_.mem_left_track_41.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_81.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__4_.mem_left_track_81.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__4_.mem_left_track_89.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__4_.mem_left_track_89.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_161.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__4_.mem_left_track_161.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_193.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__4_.mem_left_track_193.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__4_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__4_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__4_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_0.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__5_.mem_top_track_0.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_64.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__5_.mem_top_track_64.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_80.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__5_.mem_top_track_80.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__5_.mem_top_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_9.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_9.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_25.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_25.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_41.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_41.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_105.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_105.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_193.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_193.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_9__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_9.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__5_.mem_left_track_9.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_25.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_9__5_.mem_left_track_25.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_9__5_.mem_left_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__5_.mem_left_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_49.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__5_.mem_left_track_49.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__5_.mem_left_track_57.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__5_.mem_left_track_57.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_73.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__5_.mem_left_track_73.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__5_.mem_left_track_81.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__5_.mem_left_track_81.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_105.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__5_.mem_left_track_105.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_121.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__5_.mem_left_track_121.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__5_.mem_left_track_129.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__5_.mem_left_track_129.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_153.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__5_.mem_left_track_153.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_169.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__5_.mem_left_track_169.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_193.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__5_.mem_left_track_193.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__5_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_0.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__6_.mem_top_track_0.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_32.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__6_.mem_top_track_32.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__6_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_top_track_200.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_9__6_.mem_top_track_200.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_9__6_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_120.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__6_.mem_right_track_120.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__6_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_49.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_49.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_57.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_57.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_81.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_81.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_89.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_89.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_105.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_105.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_113.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_113.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_193.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_193.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__6_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_17.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_9__6_.mem_left_track_17.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_9__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_65.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__6_.mem_left_track_65.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__6_.mem_left_track_73.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__6_.mem_left_track_73.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__6_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__6_.mem_left_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__6_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_137.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__6_.mem_left_track_137.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_16.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_9__7_.mem_top_track_16.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_9__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_72.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__7_.mem_top_track_72.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__7_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_0.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_9__7_.mem_right_track_0.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_9__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_168.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__7_.mem_right_track_168.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__7_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_right_track_200.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_9__7_.mem_right_track_200.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_9__7_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_153.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__7_.mem_bottom_track_153.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__7_.mem_bottom_track_161.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__7_.mem_bottom_track_161.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__7_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_81.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__7_.mem_left_track_81.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__7_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_161.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_161.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_193.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_9__7_.mem_left_track_193.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_9__7_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__7_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__7_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_8.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__8_.mem_top_track_8.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__8_.mem_top_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__8_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_144.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__8_.mem_top_track_144.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__8_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_32.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_9__8_.mem_right_track_32.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_9__8_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_96.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__8_.mem_right_track_96.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__8_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_136.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_9__8_.mem_right_track_136.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_9__8_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_184.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__8_.mem_right_track_184.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__8_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_57.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__8_.mem_bottom_track_57.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__8_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_105.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__8_.mem_bottom_track_105.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__8_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_153.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__8_.mem_bottom_track_153.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__8_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_57.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__8_.mem_left_track_57.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__8_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__8_.mem_left_track_201.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_9__8_.mem_left_track_201.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_9__8_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__8_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_72.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__9_.mem_top_track_72.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__9_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_top_track_208.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__9_.mem_top_track_208.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__9_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_32.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__9_.mem_right_track_32.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__9_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_17.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_17.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_65.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_65.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_89.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_89.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_105.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_105.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_153.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_153.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_9__9_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_9.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__9_.mem_left_track_9.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__9_.mem_left_track_17.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_9__9_.mem_left_track_17.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_9__9_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_9__9_.mem_left_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_9__9_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_57.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_9__9_.mem_left_track_57.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_9__9_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_129.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_9__9_.mem_left_track_129.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_9__9_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__9_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__9_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_48.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_9__10_.mem_right_track_48.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_9__10_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_21.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_21.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_95.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_95.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_139.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_139.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_141.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_141.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_167.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_167.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_9__10_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_17.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_9__10_.mem_left_track_17.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_9__10_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_41.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_9__10_.mem_left_track_41.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_9__10_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_73.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_9__10_.mem_left_track_73.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_9__10_.mem_left_track_81.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_9__10_.mem_left_track_81.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_9__10_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_185.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_9__10_.mem_left_track_185.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_9__10_.mem_left_track_193.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_9__10_.mem_left_track_193.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_9__10_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_9__10_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_9__10_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_18.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_44.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_top_track_44.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_100.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_top_track_100.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_top_track_102.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_top_track_102.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_130.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_top_track_130.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_176.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_top_track_176.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_top_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_top_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_15.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_left_track_15.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_19.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_111.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_left_track_111.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_139.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_10__0_.mem_left_track_139.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_10__0_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_161.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_161.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_163.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_163.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__0_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__0_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_24.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_10__1_.mem_top_track_24.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_10__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_48.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_10__1_.mem_top_track_48.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_10__1_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_80.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__1_.mem_top_track_80.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__1_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_136.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_136.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_49.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__1_.mem_bottom_track_49.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__1_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_113.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_10__1_.mem_bottom_track_113.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_10__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_7.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_11.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_13.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_15.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_19.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_21.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_23.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_27.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__1_.mem_left_track_27.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__1_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_29.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_31.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_31.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_37.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_39.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_39.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_43.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_43.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_45.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_47.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_47.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_55.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_55.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_57.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__1_.mem_left_track_57.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__1_.mem_left_track_59.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_59.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_61.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_61.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_63.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_63.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_67.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_67.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_75.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_75.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_77.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_77.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_79.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_79.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_81.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__1_.mem_left_track_81.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__1_.mem_left_track_83.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_83.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_85.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_85.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_87.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_87.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_91.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_91.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_93.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_93.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_95.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_95.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_99.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_99.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_101.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_101.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_103.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_103.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_109.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_109.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_111.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_111.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_115.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_115.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_117.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_117.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_119.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_119.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_127.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_127.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_131.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_131.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_133.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_133.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_135.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_135.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_139.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_139.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_147.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_147.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_149.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_149.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_151.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_151.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_155.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_155.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_157.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_157.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_165.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_165.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_167.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_167.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_171.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_171.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_173.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_173.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_175.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_175.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_181.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_181.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_183.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_183.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_187.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_187.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_189.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_189.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_191.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_191.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_199.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_199.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_203.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_203.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_205.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_205.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_207.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_207.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__1_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__1_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_16.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__2_.mem_top_track_16.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_136.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_136.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_9.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_9.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_49.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_49.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_105.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_105.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_161.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_161.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_177.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_177.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__2_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_13.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__2_.mem_left_track_13.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__2_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_21.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_21.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_27.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__2_.mem_left_track_27.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__2_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_39.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_10__2_.mem_left_track_39.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_10__2_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_77.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_77.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_103.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__2_.mem_left_track_103.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__2_.mem_left_track_105.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__2_.mem_left_track_105.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__2_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_155.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_10__2_.mem_left_track_155.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_10__2_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_175.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_10__2_.mem_left_track_175.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_10__2_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_191.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_191.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__2_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__2_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_48.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__3_.mem_top_track_48.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__3_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_120.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_144.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__3_.mem_top_track_144.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__3_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_192.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__3_.mem_top_track_192.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_208.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_top_track_208.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_121.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_129.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_10__3_.mem_bottom_track_129.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_10__3_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_65.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__3_.mem_left_track_65.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__3_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_183.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_183.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__3_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__3_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_32.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_32.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_56.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__4_.mem_top_track_56.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__4_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_120.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_120.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_136.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__4_.mem_top_track_136.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__4_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_9.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__4_.mem_bottom_track_9.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_73.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__4_.mem_bottom_track_73.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__4_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_105.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__4_.mem_bottom_track_105.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__4_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_161.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_177.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_47.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__4_.mem_left_track_47.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__4_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_55.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__4_.mem_left_track_55.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__4_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_93.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__4_.mem_left_track_93.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__4_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_107.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__4_.mem_left_track_107.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__4_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_157.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_157.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_169.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__4_.mem_left_track_169.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__4_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__4_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__4_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_72.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_10__5_.mem_top_track_72.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_10__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_136.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_10__5_.mem_top_track_136.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_10__5_.mem_top_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_10__5_.mem_top_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_10__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_184.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_10__5_.mem_top_track_184.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_10__5_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_57.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__5_.mem_bottom_track_57.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__5_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_73.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_153.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__5_.mem_bottom_track_153.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__5_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_193.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__5_.mem_bottom_track_193.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__5_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_21.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_27.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_27.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_29.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_35.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_35.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_47.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_47.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_51.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_51.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_53.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_53.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_63.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_63.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_67.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_67.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_69.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_69.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_83.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_83.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_85.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_85.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_87.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_87.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_99.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_99.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_101.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_101.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_103.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_103.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_107.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_107.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_117.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_117.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_123.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_123.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_135.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_135.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_141.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_141.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_143.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_143.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_147.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_147.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_149.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_149.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_151.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_151.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_155.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_155.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_157.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_157.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_163.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_163.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_165.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_165.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_167.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_167.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_171.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_171.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_173.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_173.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_175.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_175.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_179.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_179.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_181.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_181.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_183.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_183.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_187.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_187.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_189.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_189.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_191.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_191.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_195.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_195.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_197.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_197.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_199.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_199.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_203.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_203.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_205.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_205.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_207.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_207.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__5_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__5_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_24.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_24.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_112.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_112.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_168.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__6_.mem_top_track_168.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__6_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_208.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_top_track_208.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_25.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_10__6_.mem_bottom_track_25.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_10__6_.mem_bottom_track_33.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_21.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_23.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_27.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_27.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_29.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_35.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_35.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_47.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_47.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_53.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_67.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_67.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_69.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_69.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_85.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_85.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_87.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_87.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_99.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_99.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_101.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_101.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_103.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_103.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_107.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_107.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_119.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_119.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_123.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_123.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_125.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_125.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_139.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_139.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_141.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_141.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_143.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_143.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_147.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_147.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_149.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_149.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_151.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_151.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_155.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_155.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_157.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_157.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_159.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_159.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_163.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_163.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_165.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_165.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_167.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_167.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_171.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_171.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_173.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_173.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_175.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_175.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_179.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_179.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_181.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_181.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_183.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_183.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_187.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_187.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_189.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_189.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_191.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_191.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_195.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_195.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_197.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_197.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_199.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_199.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_203.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_203.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_205.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_205.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_207.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_207.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_10__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_0.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__7_.mem_top_track_0.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__7_.mem_top_track_8.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__7_.mem_top_track_8.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__7_.mem_top_track_16.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_16.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_56.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_56.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_120.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_120.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_184.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__7_.mem_top_track_184.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__7_.mem_top_track_192.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__7_.mem_top_track_192.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__7_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_208.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_top_track_208.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_97.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_97.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_129.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_129.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_145.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_145.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_177.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_177.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_185.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_185.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__7_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_31.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_31.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_55.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__7_.mem_left_track_55.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__7_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_87.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__7_.mem_left_track_87.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__7_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__7_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__7_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_40.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_40.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_48.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_10__8_.mem_top_track_48.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_10__8_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_80.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__8_.mem_top_track_80.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__8_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_152.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_152.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_17.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_17.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_57.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_57.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_81.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_81.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_105.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_105.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_121.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_121.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__8_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_169.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_23.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_23.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_33.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__8_.mem_left_track_33.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__8_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_45.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_45.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_55.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__8_.mem_left_track_55.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__8_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_93.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__8_.mem_left_track_93.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__8_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_109.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__8_.mem_left_track_109.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__8_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_161.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__8_.mem_left_track_161.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__8_.mem_left_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__8_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__8_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_64.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_10__9_.mem_top_track_64.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_10__9_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_88.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_10__9_.mem_top_track_88.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_10__9_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_9.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_10__9_.mem_bottom_track_9.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_10__9_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_21.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__9_.mem_left_track_21.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__9_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_33.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_33.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_85.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_85.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_117.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__9_.mem_left_track_117.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__9_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_185.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__9_.mem_left_track_185.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__9_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_191.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__9_.mem_left_track_191.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__9_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_201.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_201.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__9_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__9_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_13.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_87.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_111.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_169.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__10_.mem_bottom_track_169.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__10_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_205.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_67.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_67.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_69.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__10_.mem_left_track_69.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__10_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_85.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_85.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_167.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_10__10_.mem_left_track_167.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_10__10_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_191.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_191.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_10__10_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_10__10_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_0.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_1.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_7.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_1__10_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_1__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_1__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_5.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_5.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_1.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_2.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_3.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_4.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_6.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_7.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_2__10_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_2__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_2__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_2__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_7.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_4.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_4.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_3.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_6.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_3__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_1.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_2.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_4__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_2.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_4.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_5.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_7.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_3.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_5.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_0.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_1.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_1.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_2.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_2.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_0.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_0.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_4.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_5.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_5__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_5__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_4.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_5.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_6.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_7.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_6__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_2.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_3.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_4.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_5.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_6.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_7.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_8.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_8.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_9.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_9.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_10.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_10.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_11.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_11.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_12.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_12.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_13.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_13.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_14.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_14.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_15.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_15.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_16.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_16.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_17.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_17.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_18.mem_out[0:4] = 5'b10100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_18.mem_outb[0:4] = 5'b01011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_19.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_19.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_20.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_20.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_21.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_21.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_22.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_22.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_23.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_23.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_24.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_24.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_25.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_25.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_26.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_26.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_27.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_27.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_28.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_28.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_29.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_29.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_30.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_30.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_31.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_31.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_32.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_32.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_33.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_33.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_34.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_34.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_35.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_35.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_36.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_36.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_37.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_37.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_38.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_38.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_39.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_39.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_40.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_40.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_41.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_41.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_42.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_42.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_43.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_43.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_44.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_44.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_45.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_45.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_46.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_46.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_47.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_47.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_48.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_48.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_49.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_49.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_50.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_50.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_51.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cbx_6__5_.mem_bottom_ipin_51.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_6__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_0.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_0.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_1.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_1.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_2.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_2.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_3.mem_out[0:5] = 6'b100111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_3.mem_outb[0:5] = 6'b011000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_4.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_4.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_5.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_5.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_6.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_6.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_7.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_7.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_8.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_8.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_9.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_9.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_10.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_10.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_11.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_11.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_12.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_12.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_13.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_13.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_14.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_14.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_15.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_15.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_16.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_16.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_17.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_17.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_18.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_18.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_19.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_19.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_20.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_20.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_21.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_21.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_22.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_22.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_23.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_23.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_24.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_24.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_25.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_25.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_26.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_26.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_27.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_27.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_28.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_28.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_29.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_29.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_30.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_30.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_31.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_31.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_32.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_32.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_33.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_33.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_34.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_34.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_35.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_35.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_36.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_36.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_37.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_37.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_38.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_38.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_39.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_39.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_40.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_40.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_41.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_41.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_42.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_42.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_43.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_43.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_44.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_44.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_45.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_45.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_46.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_46.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_47.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_47.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_48.mem_out[0:5] = 6'b100111;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_48.mem_outb[0:5] = 6'b011000;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_49.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_49.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_50.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_50.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_51.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_51.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_52.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_52.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_6__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_6__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_1.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_3.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_5.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_7.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cbx_6__10_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cbx_6__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_6__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_6__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_6__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_1.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_0.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_1.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_6.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_7.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_0.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_4.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_4.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_5.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_5.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_0.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_1.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_2.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_3.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_4.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__10_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_7__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_7__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_7__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_5.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_7.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_5.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_0.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_7.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_7.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cbx_8__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_0.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_0.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_2.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_6.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_8__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_8__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_0.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_1.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_2.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_6.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_7.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cbx_9__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_0.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_6.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_6.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__2_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_1.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_4.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_6.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_9__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_9__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_0.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_1.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_3.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_6.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__0_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_0.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_1.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_1.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_4.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_4.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__1_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_7.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cbx_10__2_.mem_top_ipin_7.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cbx_10__3_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__3_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__3_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__3_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__3_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__3_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__3_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__3_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__4_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__4_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__4_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__4_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__4_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__4_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__4_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__4_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_10.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_10.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_11.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_11.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_12.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_12.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_13.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_13.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_14.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_14.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_15.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_15.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_16.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_16.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_19.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_19.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_20.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_20.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_21.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_21.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_22.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_22.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_23.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_23.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_24.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_24.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_27.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_27.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_28.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_28.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_29.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_29.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_30.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_30.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_31.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_31.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_32.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_32.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_33.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_33.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_36.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_36.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_37.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_37.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_38.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_38.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_39.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_39.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_40.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_40.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_41.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_41.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_42.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_42.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_45.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_45.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_46.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_46.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_47.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_47.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_48.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_48.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_49.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_49.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_50.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_50.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_51.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_bottom_ipin_51.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_10.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_10.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_11.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_11.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_12.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_12.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_13.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_13.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_14.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_14.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_15.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_15.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_16.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_16.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_19.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_19.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_20.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_20.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_21.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_21.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_22.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_22.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_23.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_23.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_24.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_24.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_25.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_25.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_28.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_28.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_29.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_29.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_30.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_30.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_31.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_31.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_32.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_32.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_33.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_33.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_34.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_34.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_37.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_37.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_38.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_38.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_39.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_39.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_40.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_40.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_41.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_41.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_42.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_42.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_45.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_45.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_46.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_46.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_47.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_47.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_48.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_48.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_49.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_49.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_50.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_50.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_51.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_51.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_52.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__6_.mem_top_ipin_52.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__7_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__7_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__7_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__7_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__7_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__7_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__7_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__7_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__7_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__7_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__8_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__8_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__8_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__8_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__8_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__8_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__8_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__8_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__8_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__8_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__9_.mem_bottom_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__9_.mem_bottom_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__9_.mem_bottom_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__9_.mem_bottom_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__9_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__9_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__9_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__9_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__9_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__9_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_0.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_1.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_3.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_5.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_6.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__10_.mem_bottom_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__10_.mem_top_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__10_.mem_top_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__10_.mem_top_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cbx_10__10_.mem_top_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cbx_10__10_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_10__10_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cby_0__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cby_0__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_2.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_2.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_3.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_3.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_5.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_1.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_1.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_2.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_2.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_5.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_5.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_6.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_6.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cby_0__8_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_1.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cby_0__9_.mem_right_ipin_1.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cby_0__9_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_3.mem_out[0:5] = 6'b100111;
	force U0_formal_verification.cby_0__9_.mem_right_ipin_3.mem_outb[0:5] = 6'b011000;
	force U0_formal_verification.cby_0__9_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__9_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_0.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cby_0__10_.mem_right_ipin_0.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cby_0__10_.mem_right_ipin_1.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cby_0__10_.mem_right_ipin_1.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cby_0__10_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_0__10_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_6.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_1__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_1__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:5] = 6'b100100;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_2__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_2__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_6.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_6.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_3.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_3__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_3__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_7.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cby_3__1_.mem_right_ipin_7.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_3.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_3.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_5.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_5.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_3__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_3__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_3.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_4__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_4__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_4__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_4__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_0.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_5__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_5__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_left_ipin_7.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_5__1_.mem_left_ipin_7.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_4.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_4.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_6.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_6.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__6_.mem_left_ipin_0.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_0.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_1.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_1.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_2.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_2.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_3.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_3.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_4.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_4.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_5.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_5.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_6.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_6.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_7.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_7.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_8.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_8.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_9.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_9.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_10.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_10.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_11.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_11.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_12.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_12.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_13.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_13.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_14.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_14.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_15.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_15.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_16.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_16.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_17.mem_out[0:4] = 5'b11000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_17.mem_outb[0:4] = 5'b00111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_18.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_18.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_19.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_19.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_20.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_20.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_21.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_21.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_22.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_22.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_23.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_23.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_24.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_24.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_25.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_25.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_26.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_26.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_27.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_27.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_28.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_28.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_29.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_29.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_30.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_30.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_31.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_31.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_32.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_32.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_33.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_33.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_34.mem_out[0:4] = 5'b11100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_34.mem_outb[0:4] = 5'b00011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_35.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_35.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_36.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_36.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_37.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_37.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_38.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_38.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_39.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_39.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_40.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_40.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_41.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_41.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_42.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_42.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_43.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_43.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_44.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_44.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_45.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_45.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_46.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_46.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_47.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_47.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_50.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__6_.mem_left_ipin_50.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_left_ipin_51.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cby_5__6_.mem_left_ipin_51.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cby_5__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_5__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_5__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_5__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_5__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_3.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_6__1_.mem_left_ipin_3.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_6__1_.mem_left_ipin_4.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cby_6__1_.mem_left_ipin_4.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cby_6__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_6.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_6__1_.mem_left_ipin_6.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_6__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_5.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_6__1_.mem_right_ipin_5.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_6__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_3.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_3.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_6.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_5.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_5.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_6.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_6.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_0.mem_out[0:5] = 6'b000101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_0.mem_outb[0:5] = 6'b111010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_1.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_1.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_2.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_2.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_3.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_3.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_4.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_4.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_5.mem_out[0:5] = 6'b100111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_5.mem_outb[0:5] = 6'b011000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_7.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_7.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_8.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_8.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_9.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_9.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_10.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_10.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_11.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_11.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_12.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_12.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_13.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_13.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_14.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_14.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_15.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_15.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_16.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_16.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_17.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_17.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_18.mem_out[0:4] = 5'b11100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_18.mem_outb[0:4] = 5'b00011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_19.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_19.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_20.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_20.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_21.mem_out[0:5] = 6'b001000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_21.mem_outb[0:5] = 6'b110111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_22.mem_out[0:5] = 6'b100111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_22.mem_outb[0:5] = 6'b011000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_23.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_23.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_24.mem_out[0:5] = 6'b011100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_24.mem_outb[0:5] = 6'b100011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_25.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_25.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_26.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_26.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_27.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_27.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_28.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_28.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_29.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_29.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_30.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_30.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_31.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_31.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_32.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_32.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_33.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_33.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_34.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_34.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_35.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_35.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_36.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_36.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_37.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_37.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_38.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_38.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_39.mem_out[0:5] = 6'b000011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_39.mem_outb[0:5] = 6'b111100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_41.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_41.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_42.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_42.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_43.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_43.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_44.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_44.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_45.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_45.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_46.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_46.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_47.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_47.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_48.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_48.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_49.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_49.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_50.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_50.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_51.mem_out[0:5] = 6'b110111;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_51.mem_outb[0:5] = 6'b001000;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_52.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cby_6__6_.mem_right_ipin_52.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cby_6__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_6__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_6__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_6__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_6__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_0.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cby_7__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cby_7__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_7.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cby_7__1_.mem_right_ipin_7.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_1.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_1.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_6.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_7.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_7.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_7__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_7__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_7__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_7__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_1.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_1.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_2.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_2.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_3.mem_out[0:5] = 6'b010000;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_3.mem_outb[0:5] = 6'b101111;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_5.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_5.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_7.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_8__1_.mem_left_ipin_7.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_8__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_4.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_8__1_.mem_right_ipin_4.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_8__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_4.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cby_8__2_.mem_left_ipin_4.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cby_8__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_8__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_8__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_8__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_8__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_3.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_9__2_.mem_left_ipin_3.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_9__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_6.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cby_9__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cby_9__2_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_2.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cby_9__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cby_9__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__3_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__3_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__3_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__3_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__4_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__4_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__4_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__4_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__5_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__5_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_10.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_10.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_11.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_11.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_12.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_12.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_13.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_13.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_14.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_14.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_15.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_15.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_18.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_18.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_19.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_19.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_20.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_20.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_21.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_21.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_22.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_22.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_23.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_23.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_24.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_24.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_27.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_27.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_28.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_28.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_29.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_29.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_30.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_30.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_31.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_31.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_32.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_32.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_33.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_33.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_36.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_36.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_37.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_37.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_38.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_38.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_39.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_39.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_40.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_40.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_41.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_41.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_42.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_42.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_45.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_45.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_46.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_46.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_47.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_47.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_48.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_48.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_49.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_49.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_50.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_50.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_51.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_left_ipin_51.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__7_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__7_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__7_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__7_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__9_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__9_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_9__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_9__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_9__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_9__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_6.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_10__1_.mem_right_ipin_6.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_10__1_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__1_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_1.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cby_10__2_.mem_left_ipin_1.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cby_10__2_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_left_ipin_7.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cby_10__2_.mem_left_ipin_7.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cby_10__2_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_1.mem_out[0:5] = 6'b001111;
	force U0_formal_verification.cby_10__2_.mem_right_ipin_1.mem_outb[0:5] = 6'b110000;
	force U0_formal_verification.cby_10__2_.mem_right_ipin_2.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cby_10__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_10__2_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__2_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__3_.mem_left_ipin_0.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_0.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_1.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_1.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_2.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_2.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_3.mem_out[0:5] = 6'b000111;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_3.mem_outb[0:5] = 6'b111000;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_4.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_4.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_5.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_5.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_10__3_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__3_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__3_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__3_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__3_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__3_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__3_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__3_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_0.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cby_10__4_.mem_left_ipin_0.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cby_10__4_.mem_left_ipin_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cby_10__4_.mem_left_ipin_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_10__4_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_6.mem_out[0:5] = 6'b011101;
	force U0_formal_verification.cby_10__4_.mem_left_ipin_6.mem_outb[0:5] = 6'b100010;
	force U0_formal_verification.cby_10__4_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__5_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__5_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__5_.mem_left_ipin_1.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_1.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_2.mem_out[0:5] = 6'b001110;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_2.mem_outb[0:5] = 6'b110001;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__5_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__5_.mem_left_ipin_4.mem_out[0:5] = 6'b001011;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_4.mem_outb[0:5] = 6'b110100;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__5_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__5_.mem_left_ipin_6.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_6.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_7.mem_out[0:5] = 6'b010101;
	force U0_formal_verification.cby_10__5_.mem_left_ipin_7.mem_outb[0:5] = 6'b101010;
	force U0_formal_verification.cby_10__5_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__5_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__5_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__5_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_left_ipin_2.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_2.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_3.mem_out[0:5] = 6'b011000;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_3.mem_outb[0:5] = 6'b100111;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_left_ipin_5.mem_out[0:5] = 6'b010110;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_5.mem_outb[0:5] = 6'b101001;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_6.mem_out[0:5] = 6'b010011;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_6.mem_outb[0:5] = 6'b101100;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_7.mem_out[0:5] = 6'b011001;
	force U0_formal_verification.cby_10__6_.mem_left_ipin_7.mem_outb[0:5] = 6'b100110;
	force U0_formal_verification.cby_10__6_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_10.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_10.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_11.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_11.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_12.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_12.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_13.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_13.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_14.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_14.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_15.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_15.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_16.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_16.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_19.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_19.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_20.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_20.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_21.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_21.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_22.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_22.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_23.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_23.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_24.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_24.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_25.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_25.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_28.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_28.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_29.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_29.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_30.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_30.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_31.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_31.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_32.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_32.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_33.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_33.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_36.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_36.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_37.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_37.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_38.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_38.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_39.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_39.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_40.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_40.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_41.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_41.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_42.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_42.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_45.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_45.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_46.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_46.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_47.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_47.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_48.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_48.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_49.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_49.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_50.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_50.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_51.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_51.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_52.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__6_.mem_right_ipin_52.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__7_.mem_left_ipin_0.mem_out[0:5] = 6'b011010;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_0.mem_outb[0:5] = 6'b100101;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_1.mem_out[0:5] = 6'b011110;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_1.mem_outb[0:5] = 6'b100001;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__7_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__7_.mem_left_ipin_3.mem_out[0:5] = 6'b010111;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_3.mem_outb[0:5] = 6'b101000;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__7_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__7_.mem_left_ipin_5.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_5.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_6.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_6.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.cby_10__7_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__7_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__7_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__7_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__7_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__7_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__7_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__7_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_0.mem_out[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_2.mem_out[0:5] = 6'b000110;
	force U0_formal_verification.cby_10__8_.mem_left_ipin_2.mem_outb[0:5] = 6'b111001;
	force U0_formal_verification.cby_10__8_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_4.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cby_10__8_.mem_left_ipin_4.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cby_10__8_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__8_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__8_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_1.mem_out[0:5] = 6'b000100;
	force U0_formal_verification.cby_10__9_.mem_left_ipin_1.mem_outb[0:5] = 6'b111011;
	force U0_formal_verification.cby_10__9_.mem_left_ipin_2.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_2.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__9_.mem_left_ipin_5.mem_out[0:5] = 6'b101111;
	force U0_formal_verification.cby_10__9_.mem_left_ipin_5.mem_outb[0:5] = 6'b010000;
	force U0_formal_verification.cby_10__9_.mem_left_ipin_6.mem_out[0:5] = 6'b111011;
	force U0_formal_verification.cby_10__9_.mem_left_ipin_6.mem_outb[0:5] = 6'b000100;
	force U0_formal_verification.cby_10__9_.mem_left_ipin_7.mem_out[0:5] = 6'b011111;
	force U0_formal_verification.cby_10__9_.mem_left_ipin_7.mem_outb[0:5] = 6'b100000;
	force U0_formal_verification.cby_10__9_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__9_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__9_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__9_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__9_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__9_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_2.mem_out[0:5] = 6'b001101;
	force U0_formal_verification.cby_10__10_.mem_left_ipin_2.mem_outb[0:5] = 6'b110010;
	force U0_formal_verification.cby_10__10_.mem_left_ipin_3.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_3.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_4.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_4.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_5.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_5.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_6.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_6.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_7.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_left_ipin_7.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_right_ipin_0.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_right_ipin_0.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_right_ipin_1.mem_out[0:5] = {6{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_right_ipin_1.mem_outb[0:5] = {6{1'b1}};
	force U0_formal_verification.cby_10__10_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_10__10_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
end
// ----- End assign bitstream to configuration memories -----
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for router_bench_top_formal_verification -----

//----- Default net type -----
`default_nettype wire

