//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[18][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul 21 20:26:54 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_18__0_ -----
module sb_18__0_(prog_clk,
                 chany_top_in,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                 chanx_left_in,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                 ccff_head,
                 chany_top_out,
                 chanx_left_out,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:105] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:105] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:105] chany_top_out;
//----- OUTPUT PORTS -----
output [0:105] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_16_sram;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_17_sram;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_18_sram;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_19_sram;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_20_sram;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_21_sram;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_22_sram;
wire [0:1] mux_tree_tapbuf_size2_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_23_sram;
wire [0:1] mux_tree_tapbuf_size2_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_24_sram;
wire [0:1] mux_tree_tapbuf_size2_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_25_sram;
wire [0:1] mux_tree_tapbuf_size2_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_26_sram;
wire [0:1] mux_tree_tapbuf_size2_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_27_sram;
wire [0:1] mux_tree_tapbuf_size2_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_28_sram;
wire [0:1] mux_tree_tapbuf_size2_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_29_sram;
wire [0:1] mux_tree_tapbuf_size2_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_30_sram;
wire [0:1] mux_tree_tapbuf_size2_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_31_sram;
wire [0:1] mux_tree_tapbuf_size2_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_32_sram;
wire [0:1] mux_tree_tapbuf_size2_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_33_sram;
wire [0:1] mux_tree_tapbuf_size2_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_34_sram;
wire [0:1] mux_tree_tapbuf_size2_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_35_sram;
wire [0:1] mux_tree_tapbuf_size2_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_36_sram;
wire [0:1] mux_tree_tapbuf_size2_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_37_sram;
wire [0:1] mux_tree_tapbuf_size2_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_38_sram;
wire [0:1] mux_tree_tapbuf_size2_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_39_sram;
wire [0:1] mux_tree_tapbuf_size2_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_100_sram;
wire [0:1] mux_tree_tapbuf_size3_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_101_sram;
wire [0:1] mux_tree_tapbuf_size3_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_102_sram;
wire [0:1] mux_tree_tapbuf_size3_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_103_sram;
wire [0:1] mux_tree_tapbuf_size3_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_104_sram;
wire [0:1] mux_tree_tapbuf_size3_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_105_sram;
wire [0:1] mux_tree_tapbuf_size3_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_106_sram;
wire [0:1] mux_tree_tapbuf_size3_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_107_sram;
wire [0:1] mux_tree_tapbuf_size3_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_108_sram;
wire [0:1] mux_tree_tapbuf_size3_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_109_sram;
wire [0:1] mux_tree_tapbuf_size3_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_110_sram;
wire [0:1] mux_tree_tapbuf_size3_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_111_sram;
wire [0:1] mux_tree_tapbuf_size3_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_112_sram;
wire [0:1] mux_tree_tapbuf_size3_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_113_sram;
wire [0:1] mux_tree_tapbuf_size3_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_114_sram;
wire [0:1] mux_tree_tapbuf_size3_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_115_sram;
wire [0:1] mux_tree_tapbuf_size3_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_116_sram;
wire [0:1] mux_tree_tapbuf_size3_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_117_sram;
wire [0:1] mux_tree_tapbuf_size3_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_118_sram;
wire [0:1] mux_tree_tapbuf_size3_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_119_sram;
wire [0:1] mux_tree_tapbuf_size3_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_120_sram;
wire [0:1] mux_tree_tapbuf_size3_120_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_121_sram;
wire [0:1] mux_tree_tapbuf_size3_121_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_122_sram;
wire [0:1] mux_tree_tapbuf_size3_122_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_123_sram;
wire [0:1] mux_tree_tapbuf_size3_123_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_124_sram;
wire [0:1] mux_tree_tapbuf_size3_124_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_125_sram;
wire [0:1] mux_tree_tapbuf_size3_125_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_126_sram;
wire [0:1] mux_tree_tapbuf_size3_126_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_127_sram;
wire [0:1] mux_tree_tapbuf_size3_127_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_128_sram;
wire [0:1] mux_tree_tapbuf_size3_128_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_129_sram;
wire [0:1] mux_tree_tapbuf_size3_129_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_130_sram;
wire [0:1] mux_tree_tapbuf_size3_130_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_131_sram;
wire [0:1] mux_tree_tapbuf_size3_131_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_132_sram;
wire [0:1] mux_tree_tapbuf_size3_132_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_133_sram;
wire [0:1] mux_tree_tapbuf_size3_133_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_134_sram;
wire [0:1] mux_tree_tapbuf_size3_134_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_135_sram;
wire [0:1] mux_tree_tapbuf_size3_135_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_136_sram;
wire [0:1] mux_tree_tapbuf_size3_136_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_137_sram;
wire [0:1] mux_tree_tapbuf_size3_137_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_138_sram;
wire [0:1] mux_tree_tapbuf_size3_138_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_139_sram;
wire [0:1] mux_tree_tapbuf_size3_139_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_140_sram;
wire [0:1] mux_tree_tapbuf_size3_140_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_141_sram;
wire [0:1] mux_tree_tapbuf_size3_141_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_142_sram;
wire [0:1] mux_tree_tapbuf_size3_142_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_143_sram;
wire [0:1] mux_tree_tapbuf_size3_143_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_144_sram;
wire [0:1] mux_tree_tapbuf_size3_144_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_145_sram;
wire [0:1] mux_tree_tapbuf_size3_145_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_146_sram;
wire [0:1] mux_tree_tapbuf_size3_146_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_147_sram;
wire [0:1] mux_tree_tapbuf_size3_147_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_148_sram;
wire [0:1] mux_tree_tapbuf_size3_148_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_149_sram;
wire [0:1] mux_tree_tapbuf_size3_149_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_150_sram;
wire [0:1] mux_tree_tapbuf_size3_150_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_151_sram;
wire [0:1] mux_tree_tapbuf_size3_151_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_152_sram;
wire [0:1] mux_tree_tapbuf_size3_152_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_153_sram;
wire [0:1] mux_tree_tapbuf_size3_153_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_154_sram;
wire [0:1] mux_tree_tapbuf_size3_154_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_155_sram;
wire [0:1] mux_tree_tapbuf_size3_155_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_156_sram;
wire [0:1] mux_tree_tapbuf_size3_156_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_157_sram;
wire [0:1] mux_tree_tapbuf_size3_157_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_158_sram;
wire [0:1] mux_tree_tapbuf_size3_158_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_159_sram;
wire [0:1] mux_tree_tapbuf_size3_159_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_160_sram;
wire [0:1] mux_tree_tapbuf_size3_160_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_161_sram;
wire [0:1] mux_tree_tapbuf_size3_161_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_162_sram;
wire [0:1] mux_tree_tapbuf_size3_162_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_163_sram;
wire [0:1] mux_tree_tapbuf_size3_163_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_164_sram;
wire [0:1] mux_tree_tapbuf_size3_164_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_165_sram;
wire [0:1] mux_tree_tapbuf_size3_165_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_166_sram;
wire [0:1] mux_tree_tapbuf_size3_166_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_167_sram;
wire [0:1] mux_tree_tapbuf_size3_167_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_168_sram;
wire [0:1] mux_tree_tapbuf_size3_168_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_169_sram;
wire [0:1] mux_tree_tapbuf_size3_169_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_170_sram;
wire [0:1] mux_tree_tapbuf_size3_170_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_171_sram;
wire [0:1] mux_tree_tapbuf_size3_171_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_33_sram;
wire [0:1] mux_tree_tapbuf_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_34_sram;
wire [0:1] mux_tree_tapbuf_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_35_sram;
wire [0:1] mux_tree_tapbuf_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_36_sram;
wire [0:1] mux_tree_tapbuf_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_37_sram;
wire [0:1] mux_tree_tapbuf_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_38_sram;
wire [0:1] mux_tree_tapbuf_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_39_sram;
wire [0:1] mux_tree_tapbuf_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_40_sram;
wire [0:1] mux_tree_tapbuf_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_41_sram;
wire [0:1] mux_tree_tapbuf_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_42_sram;
wire [0:1] mux_tree_tapbuf_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_43_sram;
wire [0:1] mux_tree_tapbuf_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_44_sram;
wire [0:1] mux_tree_tapbuf_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_45_sram;
wire [0:1] mux_tree_tapbuf_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_46_sram;
wire [0:1] mux_tree_tapbuf_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_47_sram;
wire [0:1] mux_tree_tapbuf_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_48_sram;
wire [0:1] mux_tree_tapbuf_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_49_sram;
wire [0:1] mux_tree_tapbuf_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_50_sram;
wire [0:1] mux_tree_tapbuf_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_51_sram;
wire [0:1] mux_tree_tapbuf_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_52_sram;
wire [0:1] mux_tree_tapbuf_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_53_sram;
wire [0:1] mux_tree_tapbuf_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_54_sram;
wire [0:1] mux_tree_tapbuf_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_55_sram;
wire [0:1] mux_tree_tapbuf_size3_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_56_sram;
wire [0:1] mux_tree_tapbuf_size3_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_57_sram;
wire [0:1] mux_tree_tapbuf_size3_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_58_sram;
wire [0:1] mux_tree_tapbuf_size3_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_59_sram;
wire [0:1] mux_tree_tapbuf_size3_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_60_sram;
wire [0:1] mux_tree_tapbuf_size3_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_61_sram;
wire [0:1] mux_tree_tapbuf_size3_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_62_sram;
wire [0:1] mux_tree_tapbuf_size3_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_63_sram;
wire [0:1] mux_tree_tapbuf_size3_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_64_sram;
wire [0:1] mux_tree_tapbuf_size3_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_65_sram;
wire [0:1] mux_tree_tapbuf_size3_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_66_sram;
wire [0:1] mux_tree_tapbuf_size3_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_67_sram;
wire [0:1] mux_tree_tapbuf_size3_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_68_sram;
wire [0:1] mux_tree_tapbuf_size3_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_69_sram;
wire [0:1] mux_tree_tapbuf_size3_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_70_sram;
wire [0:1] mux_tree_tapbuf_size3_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_71_sram;
wire [0:1] mux_tree_tapbuf_size3_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_72_sram;
wire [0:1] mux_tree_tapbuf_size3_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_73_sram;
wire [0:1] mux_tree_tapbuf_size3_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_74_sram;
wire [0:1] mux_tree_tapbuf_size3_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_75_sram;
wire [0:1] mux_tree_tapbuf_size3_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_76_sram;
wire [0:1] mux_tree_tapbuf_size3_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_77_sram;
wire [0:1] mux_tree_tapbuf_size3_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_78_sram;
wire [0:1] mux_tree_tapbuf_size3_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_79_sram;
wire [0:1] mux_tree_tapbuf_size3_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_80_sram;
wire [0:1] mux_tree_tapbuf_size3_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_81_sram;
wire [0:1] mux_tree_tapbuf_size3_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_82_sram;
wire [0:1] mux_tree_tapbuf_size3_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_83_sram;
wire [0:1] mux_tree_tapbuf_size3_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_84_sram;
wire [0:1] mux_tree_tapbuf_size3_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_85_sram;
wire [0:1] mux_tree_tapbuf_size3_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_86_sram;
wire [0:1] mux_tree_tapbuf_size3_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_87_sram;
wire [0:1] mux_tree_tapbuf_size3_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_88_sram;
wire [0:1] mux_tree_tapbuf_size3_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_89_sram;
wire [0:1] mux_tree_tapbuf_size3_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_90_sram;
wire [0:1] mux_tree_tapbuf_size3_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_91_sram;
wire [0:1] mux_tree_tapbuf_size3_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_92_sram;
wire [0:1] mux_tree_tapbuf_size3_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_93_sram;
wire [0:1] mux_tree_tapbuf_size3_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_94_sram;
wire [0:1] mux_tree_tapbuf_size3_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_95_sram;
wire [0:1] mux_tree_tapbuf_size3_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_96_sram;
wire [0:1] mux_tree_tapbuf_size3_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_97_sram;
wire [0:1] mux_tree_tapbuf_size3_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_98_sram;
wire [0:1] mux_tree_tapbuf_size3_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_99_sram;
wire [0:1] mux_tree_tapbuf_size3_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_136_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_137_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_138_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_139_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_140_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_141_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_142_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_143_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_144_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_145_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_146_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_147_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_148_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_149_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_150_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_151_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_152_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_153_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_154_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_155_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_156_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_157_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_158_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_159_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_160_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_161_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_162_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_163_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_164_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_165_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_166_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_167_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_168_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_169_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_170_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size3 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[0]}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size3 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[105]}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_size3 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_size3 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_size3 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size3 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_size3 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_size3 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_size3 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size3 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[97]}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_size3 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[96]}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_size3 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_size3 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size3 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_size3 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_size3 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_size3 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_size3 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_size3 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size3 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_tree_tapbuf_size3 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_tree_tapbuf_size3 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_size3 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size3 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_size3 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size3 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_tree_tapbuf_size3 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_tree_tapbuf_size3 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_size3 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size3 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_tree_tapbuf_size3 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size3 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_tree_tapbuf_size3 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chany_top_out[38]));

	mux_tree_tapbuf_size3 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_33_sram_inv[0:1]),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_size3 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_34_sram_inv[0:1]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size3 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_35_sram_inv[0:1]),
		.out(chany_top_out[41]));

	mux_tree_tapbuf_size3 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_36_sram_inv[0:1]),
		.out(chany_top_out[42]));

	mux_tree_tapbuf_size3 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_37_sram_inv[0:1]),
		.out(chany_top_out[45]));

	mux_tree_tapbuf_size3 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_38_sram_inv[0:1]),
		.out(chany_top_out[46]));

	mux_tree_tapbuf_size3 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_39_sram_inv[0:1]),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_size3 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_40_sram_inv[0:1]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size3 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_41_sram_inv[0:1]),
		.out(chany_top_out[49]));

	mux_tree_tapbuf_size3 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_42_sram_inv[0:1]),
		.out(chany_top_out[50]));

	mux_tree_tapbuf_size3 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_43_sram_inv[0:1]),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_size3 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_44_sram_inv[0:1]),
		.out(chany_top_out[54]));

	mux_tree_tapbuf_size3 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_45_sram_inv[0:1]),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_size3 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_46_sram_inv[0:1]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size3 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_47_sram_inv[0:1]),
		.out(chany_top_out[57]));

	mux_tree_tapbuf_size3 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_48_sram_inv[0:1]),
		.out(chany_top_out[58]));

	mux_tree_tapbuf_size3 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_49_sram_inv[0:1]),
		.out(chany_top_out[59]));

	mux_tree_tapbuf_size3 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_50_sram_inv[0:1]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size3 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_51_sram_inv[0:1]),
		.out(chany_top_out[63]));

	mux_tree_tapbuf_size3 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_52_sram_inv[0:1]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size3 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_53_sram_inv[0:1]),
		.out(chany_top_out[65]));

	mux_tree_tapbuf_size3 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_54_sram_inv[0:1]),
		.out(chany_top_out[66]));

	mux_tree_tapbuf_size3 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_55_sram_inv[0:1]),
		.out(chany_top_out[67]));

	mux_tree_tapbuf_size3 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_56_sram_inv[0:1]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size3 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_57_sram_inv[0:1]),
		.out(chany_top_out[69]));

	mux_tree_tapbuf_size3 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[34]}),
		.sram(mux_tree_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_58_sram_inv[0:1]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size3 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[33]}),
		.sram(mux_tree_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_59_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_tree_tapbuf_size3 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[32]}),
		.sram(mux_tree_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_60_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_tree_tapbuf_size3 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_61_sram_inv[0:1]),
		.out(chany_top_out[75]));

	mux_tree_tapbuf_size3 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[30]}),
		.sram(mux_tree_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_62_sram_inv[0:1]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size3 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[29]}),
		.sram(mux_tree_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_63_sram_inv[0:1]),
		.out(chany_top_out[77]));

	mux_tree_tapbuf_size3 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[28]}),
		.sram(mux_tree_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_64_sram_inv[0:1]),
		.out(chany_top_out[78]));

	mux_tree_tapbuf_size3 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[25]}),
		.sram(mux_tree_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_65_sram_inv[0:1]),
		.out(chany_top_out[81]));

	mux_tree_tapbuf_size3 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[24]}),
		.sram(mux_tree_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_66_sram_inv[0:1]),
		.out(chany_top_out[82]));

	mux_tree_tapbuf_size3 mux_top_track_166 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_67_sram_inv[0:1]),
		.out(chany_top_out[83]));

	mux_tree_tapbuf_size3 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[22]}),
		.sram(mux_tree_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_68_sram_inv[0:1]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size3 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[21]}),
		.sram(mux_tree_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_69_sram_inv[0:1]),
		.out(chany_top_out[85]));

	mux_tree_tapbuf_size3 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[20]}),
		.sram(mux_tree_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_70_sram_inv[0:1]),
		.out(chany_top_out[86]));

	mux_tree_tapbuf_size3 mux_top_track_174 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_71_sram_inv[0:1]),
		.out(chany_top_out[87]));

	mux_tree_tapbuf_size3 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[16]}),
		.sram(mux_tree_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_72_sram_inv[0:1]),
		.out(chany_top_out[90]));

	mux_tree_tapbuf_size3 mux_top_track_182 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_73_sram_inv[0:1]),
		.out(chany_top_out[91]));

	mux_tree_tapbuf_size3 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[14]}),
		.sram(mux_tree_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_74_sram_inv[0:1]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size3 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[13]}),
		.sram(mux_tree_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_75_sram_inv[0:1]),
		.out(chany_top_out[93]));

	mux_tree_tapbuf_size3 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[12]}),
		.sram(mux_tree_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_76_sram_inv[0:1]),
		.out(chany_top_out[94]));

	mux_tree_tapbuf_size3 mux_top_track_190 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_77_sram_inv[0:1]),
		.out(chany_top_out[95]));

	mux_tree_tapbuf_size3 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[10]}),
		.sram(mux_tree_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_78_sram_inv[0:1]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size3 mux_top_track_198 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_79_sram_inv[0:1]),
		.out(chany_top_out[99]));

	mux_tree_tapbuf_size3 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[6]}),
		.sram(mux_tree_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_80_sram_inv[0:1]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size3 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[5]}),
		.sram(mux_tree_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_81_sram_inv[0:1]),
		.out(chany_top_out[101]));

	mux_tree_tapbuf_size3 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[4]}),
		.sram(mux_tree_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_82_sram_inv[0:1]),
		.out(chany_top_out[102]));

	mux_tree_tapbuf_size3 mux_top_track_206 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_83_sram_inv[0:1]),
		.out(chany_top_out[103]));

	mux_tree_tapbuf_size3 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[2]}),
		.sram(mux_tree_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_84_sram_inv[0:1]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size3 mux_top_track_210 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[1]}),
		.sram(mux_tree_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_85_sram_inv[0:1]),
		.out(chany_top_out[105]));

	mux_tree_tapbuf_size3 mux_left_track_1 (
		.in({chany_top_in[0], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_86_sram_inv[0:1]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size3 mux_left_track_3 (
		.in({chany_top_in[105], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_87_sram_inv[0:1]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_size3 mux_left_track_5 (
		.in({chany_top_in[104], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_88_sram_inv[0:1]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_size3 mux_left_track_7 (
		.in({chany_top_in[103], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_89_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_size3 mux_left_track_9 (
		.in({chany_top_in[102], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_90_sram_inv[0:1]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size3 mux_left_track_11 (
		.in({chany_top_in[101], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_91_sram_inv[0:1]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_size3 mux_left_track_13 (
		.in({chany_top_in[100], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_92_sram_inv[0:1]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_size3 mux_left_track_15 (
		.in({chany_top_in[99], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_93_sram_inv[0:1]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_size3 mux_left_track_17 (
		.in({chany_top_in[98], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_94_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size3 mux_left_track_19 (
		.in({chany_top_in[97], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_95_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_size3 mux_left_track_21 (
		.in({chany_top_in[96], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_96_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_size3 mux_left_track_23 (
		.in({chany_top_in[95], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_97_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_size3 mux_left_track_25 (
		.in({chany_top_in[94], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_98_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size3 mux_left_track_27 (
		.in({chany_top_in[93], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_99_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_size3 mux_left_track_29 (
		.in({chany_top_in[92], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_100_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_size3 mux_left_track_31 (
		.in({chany_top_in[91], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_101_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_size3 mux_left_track_37 (
		.in({chany_top_in[88], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_102_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_size3 mux_left_track_39 (
		.in({chany_top_in[87], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_103_sram_inv[0:1]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_size3 mux_left_track_41 (
		.in({chany_top_in[86], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_104_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size3 mux_left_track_43 (
		.in({chany_top_in[85], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_105_sram_inv[0:1]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_size3 mux_left_track_45 (
		.in({chany_top_in[84], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_106_sram_inv[0:1]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_size3 mux_left_track_47 (
		.in({chany_top_in[83], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_107_sram_inv[0:1]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_size3 mux_left_track_49 (
		.in({chany_top_in[82], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_108_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size3 mux_left_track_55 (
		.in({chany_top_in[79], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_109_sram_inv[0:1]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_size3 mux_left_track_57 (
		.in({chany_top_in[78], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_110_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size3 mux_left_track_59 (
		.in({chany_top_in[77], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_111_sram_inv[0:1]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_size3 mux_left_track_61 (
		.in({chany_top_in[76], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_112_sram_inv[0:1]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_size3 mux_left_track_63 (
		.in({chany_top_in[75], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_113_sram_inv[0:1]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_size3 mux_left_track_65 (
		.in({chany_top_in[74], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_114_sram_inv[0:1]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size3 mux_left_track_67 (
		.in({chany_top_in[73], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_115_sram_inv[0:1]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_size3 mux_left_track_73 (
		.in({chany_top_in[70], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_116_sram_inv[0:1]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size3 mux_left_track_75 (
		.in({chany_top_in[69], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_117_sram_inv[0:1]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_size3 mux_left_track_77 (
		.in({chany_top_in[68], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_118_sram_inv[0:1]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_size3 mux_left_track_79 (
		.in({chany_top_in[67], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_119_sram_inv[0:1]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_size3 mux_left_track_81 (
		.in({chany_top_in[66], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_120_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_120_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size3 mux_left_track_83 (
		.in({chany_top_in[65], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_121_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_121_sram_inv[0:1]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_size3 mux_left_track_85 (
		.in({chany_top_in[64], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_122_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_122_sram_inv[0:1]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_size3 mux_left_track_91 (
		.in({chany_top_in[61], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_123_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_123_sram_inv[0:1]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_size3 mux_left_track_93 (
		.in({chany_top_in[60], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_124_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_124_sram_inv[0:1]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_size3 mux_left_track_95 (
		.in({chany_top_in[59], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_125_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_125_sram_inv[0:1]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_size3 mux_left_track_97 (
		.in({chany_top_in[58], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_126_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_126_sram_inv[0:1]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size3 mux_left_track_99 (
		.in({chany_top_in[57], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_127_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_127_sram_inv[0:1]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_size3 mux_left_track_101 (
		.in({chany_top_in[56], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_128_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_128_sram_inv[0:1]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_size3 mux_left_track_103 (
		.in({chany_top_in[55], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_129_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_129_sram_inv[0:1]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_size3 mux_left_track_109 (
		.in({chany_top_in[52], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_130_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_130_sram_inv[0:1]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_size3 mux_left_track_111 (
		.in({chany_top_in[51], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_131_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_131_sram_inv[0:1]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_size3 mux_left_track_113 (
		.in({chany_top_in[50], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_132_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_132_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size3 mux_left_track_115 (
		.in({chany_top_in[49], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_133_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_133_sram_inv[0:1]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_size3 mux_left_track_117 (
		.in({chany_top_in[48], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_134_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_134_sram_inv[0:1]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_size3 mux_left_track_119 (
		.in({chany_top_in[47], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_135_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_135_sram_inv[0:1]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_size3 mux_left_track_121 (
		.in({chany_top_in[46], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_136_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_136_sram_inv[0:1]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size3 mux_left_track_127 (
		.in({chany_top_in[43], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_137_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_137_sram_inv[0:1]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_size3 mux_left_track_129 (
		.in({chany_top_in[42], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_138_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_138_sram_inv[0:1]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size3 mux_left_track_131 (
		.in({chany_top_in[41], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_139_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_139_sram_inv[0:1]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_size3 mux_left_track_133 (
		.in({chany_top_in[40], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_140_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_140_sram_inv[0:1]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_size3 mux_left_track_135 (
		.in({chany_top_in[39], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_141_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_141_sram_inv[0:1]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_size3 mux_left_track_137 (
		.in({chany_top_in[38], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_142_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_142_sram_inv[0:1]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size3 mux_left_track_139 (
		.in({chany_top_in[37], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_143_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_143_sram_inv[0:1]),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_size3 mux_left_track_145 (
		.in({chany_top_in[34], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_144_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_144_sram_inv[0:1]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size3 mux_left_track_147 (
		.in({chany_top_in[33], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_145_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_145_sram_inv[0:1]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_size3 mux_left_track_149 (
		.in({chany_top_in[32], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_146_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_146_sram_inv[0:1]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_size3 mux_left_track_151 (
		.in({chany_top_in[31], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_147_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_147_sram_inv[0:1]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_size3 mux_left_track_153 (
		.in({chany_top_in[30], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_148_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_148_sram_inv[0:1]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size3 mux_left_track_155 (
		.in({chany_top_in[29], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_149_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_149_sram_inv[0:1]),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_size3 mux_left_track_157 (
		.in({chany_top_in[28], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_150_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_150_sram_inv[0:1]),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_size3 mux_left_track_163 (
		.in({chany_top_in[25], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_151_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_151_sram_inv[0:1]),
		.out(chanx_left_out[81]));

	mux_tree_tapbuf_size3 mux_left_track_165 (
		.in({chany_top_in[24], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_152_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_152_sram_inv[0:1]),
		.out(chanx_left_out[82]));

	mux_tree_tapbuf_size3 mux_left_track_167 (
		.in({chany_top_in[23], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_153_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_153_sram_inv[0:1]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_size3 mux_left_track_169 (
		.in({chany_top_in[22], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_154_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_154_sram_inv[0:1]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size3 mux_left_track_171 (
		.in({chany_top_in[21], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_155_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_155_sram_inv[0:1]),
		.out(chanx_left_out[85]));

	mux_tree_tapbuf_size3 mux_left_track_173 (
		.in({chany_top_in[20], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_156_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_156_sram_inv[0:1]),
		.out(chanx_left_out[86]));

	mux_tree_tapbuf_size3 mux_left_track_175 (
		.in({chany_top_in[19], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_157_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_157_sram_inv[0:1]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_size3 mux_left_track_181 (
		.in({chany_top_in[16], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_158_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_158_sram_inv[0:1]),
		.out(chanx_left_out[90]));

	mux_tree_tapbuf_size3 mux_left_track_183 (
		.in({chany_top_in[15], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_159_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_159_sram_inv[0:1]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_size3 mux_left_track_185 (
		.in({chany_top_in[14], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_160_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_160_sram_inv[0:1]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size3 mux_left_track_187 (
		.in({chany_top_in[13], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_161_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_161_sram_inv[0:1]),
		.out(chanx_left_out[93]));

	mux_tree_tapbuf_size3 mux_left_track_189 (
		.in({chany_top_in[12], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_162_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_162_sram_inv[0:1]),
		.out(chanx_left_out[94]));

	mux_tree_tapbuf_size3 mux_left_track_191 (
		.in({chany_top_in[11], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_163_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_163_sram_inv[0:1]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_size3 mux_left_track_193 (
		.in({chany_top_in[10], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_164_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_164_sram_inv[0:1]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size3 mux_left_track_199 (
		.in({chany_top_in[7], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_165_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_165_sram_inv[0:1]),
		.out(chanx_left_out[99]));

	mux_tree_tapbuf_size3 mux_left_track_201 (
		.in({chany_top_in[6], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_166_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_166_sram_inv[0:1]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size3 mux_left_track_203 (
		.in({chany_top_in[5], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_167_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_167_sram_inv[0:1]),
		.out(chanx_left_out[101]));

	mux_tree_tapbuf_size3 mux_left_track_205 (
		.in({chany_top_in[4], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_168_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_168_sram_inv[0:1]),
		.out(chanx_left_out[102]));

	mux_tree_tapbuf_size3 mux_left_track_207 (
		.in({chany_top_in[3], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_169_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_169_sram_inv[0:1]),
		.out(chanx_left_out[103]));

	mux_tree_tapbuf_size3 mux_left_track_209 (
		.in({chany_top_in[2], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_170_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_170_sram_inv[0:1]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size3 mux_left_track_211 (
		.in({chany_top_in[1], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_171_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_171_sram_inv[0:1]),
		.out(chanx_left_out[105]));

	mux_tree_tapbuf_size3_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_55_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_56_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_57_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_58_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_59_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_60_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_61_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_62_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_63_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_64_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_65_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_66_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_67_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_68_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_69_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_70_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_71_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_72_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_73_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_74_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_75_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_76_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_77_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_78_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_79_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_80_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_81_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_82_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_83_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_84_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_85_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_86_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_87_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_88_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_89_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_90_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_91_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_92_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_93_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_94_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_95_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_96_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_97_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_98_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_99_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_100_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_101_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_102_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_103_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_104_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_105_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_106_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_107_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_108_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_109_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_110_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_111_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_112_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_113_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_114_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_115_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_116_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_117_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_118_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_119_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_120_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_120_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_121_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_121_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_122_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_122_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_123_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_123_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_124_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_124_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_125_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_125_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_126_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_126_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_127_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_127_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_128_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_128_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_129_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_129_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_130_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_130_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_131_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_131_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_132_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_132_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_133_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_133_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_134_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_134_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_135_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_135_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_136_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_136_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_136_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_137_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_137_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_137_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_137_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_138_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_138_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_138_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_138_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_139_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_139_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_139_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_139_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_140_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_140_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_140_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_140_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_141_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_141_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_141_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_141_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_142_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_142_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_142_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_142_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_143_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_143_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_143_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_144_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_144_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_144_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_147 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_144_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_145_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_145_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_145_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_149 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_145_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_146_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_146_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_146_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_151 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_146_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_147_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_147_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_147_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_147_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_148_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_148_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_148_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_155 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_148_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_149_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_149_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_149_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_157 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_149_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_150_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_150_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_150_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_163 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_151_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_151_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_151_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_165 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_151_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_152_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_152_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_152_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_167 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_152_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_153_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_153_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_153_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_153_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_154_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_154_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_154_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_171 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_154_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_155_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_155_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_155_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_173 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_155_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_156_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_156_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_156_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_175 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_156_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_157_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_157_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_157_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_181 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_158_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_158_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_158_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_183 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_158_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_159_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_159_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_159_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_159_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_160_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_160_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_160_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_187 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_160_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_161_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_161_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_161_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_189 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_161_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_162_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_162_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_162_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_191 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_162_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_163_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_163_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_163_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_163_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_164_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_164_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_164_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_199 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_165_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_165_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_165_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_165_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_166_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_166_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_166_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_203 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_166_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_167_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_167_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_167_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_205 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_167_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_168_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_168_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_168_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_207 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_168_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_169_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_169_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_169_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_169_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_170_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_170_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_170_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_211 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_170_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_171_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_171_sram_inv[0:1]));

	mux_tree_tapbuf_size2 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size2 mux_top_track_34 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_size2 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_tree_tapbuf_size2 mux_top_track_52 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(chany_top_out[26]));

	mux_tree_tapbuf_size2 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_tree_tapbuf_size2 mux_top_track_70 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_size2 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_size2 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size2 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size2 mux_top_track_106 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_top_out[53]));

	mux_tree_tapbuf_size2 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_top_out[61]));

	mux_tree_tapbuf_size2 mux_top_track_124 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_top_out[62]));

	mux_tree_tapbuf_size2 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[36]}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_top_out[70]));

	mux_tree_tapbuf_size2 mux_top_track_142 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_top_out[71]));

	mux_tree_tapbuf_size2 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_tree_tapbuf_size2 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[26]}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size2 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[18]}),
		.sram(mux_tree_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size2 mux_top_track_178 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[17]}),
		.sram(mux_tree_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_top_out[89]));

	mux_tree_tapbuf_size2 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[9]}),
		.sram(mux_tree_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_18_sram_inv[0:1]),
		.out(chany_top_out[97]));

	mux_tree_tapbuf_size2 mux_top_track_196 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[8]}),
		.sram(mux_tree_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_19_sram_inv[0:1]),
		.out(chany_top_out[98]));

	mux_tree_tapbuf_size2 mux_left_track_33 (
		.in({chany_top_in[90], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_20_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size2 mux_left_track_35 (
		.in({chany_top_in[89], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_21_sram_inv[0:1]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_size2 mux_left_track_51 (
		.in({chany_top_in[81], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_22_sram_inv[0:1]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_size2 mux_left_track_53 (
		.in({chany_top_in[80], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_23_sram_inv[0:1]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_size2 mux_left_track_69 (
		.in({chany_top_in[72], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_24_sram_inv[0:1]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_size2 mux_left_track_71 (
		.in({chany_top_in[71], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_25_sram_inv[0:1]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_size2 mux_left_track_87 (
		.in({chany_top_in[63], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_26_sram_inv[0:1]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_size2 mux_left_track_89 (
		.in({chany_top_in[62], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_27_sram_inv[0:1]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size2 mux_left_track_105 (
		.in({chany_top_in[54], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_28_sram_inv[0:1]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size2 mux_left_track_107 (
		.in({chany_top_in[53], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_29_sram_inv[0:1]),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_size2 mux_left_track_123 (
		.in({chany_top_in[45], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_30_sram_inv[0:1]),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_size2 mux_left_track_125 (
		.in({chany_top_in[44], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_31_sram_inv[0:1]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_size2 mux_left_track_141 (
		.in({chany_top_in[36], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_32_sram_inv[0:1]),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_size2 mux_left_track_143 (
		.in({chany_top_in[35], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_33_sram_inv[0:1]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_size2 mux_left_track_159 (
		.in({chany_top_in[27], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_34_sram_inv[0:1]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_size2 mux_left_track_161 (
		.in({chany_top_in[26], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_35_sram_inv[0:1]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size2 mux_left_track_177 (
		.in({chany_top_in[18], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_36_sram_inv[0:1]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size2 mux_left_track_179 (
		.in({chany_top_in[17], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_37_sram_inv[0:1]),
		.out(chanx_left_out[89]));

	mux_tree_tapbuf_size2 mux_left_track_195 (
		.in({chany_top_in[9], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_38_sram_inv[0:1]),
		.out(chanx_left_out[97]));

	mux_tree_tapbuf_size2 mux_left_track_197 (
		.in({chany_top_in[8], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_39_sram_inv[0:1]),
		.out(chanx_left_out[98]));

	mux_tree_tapbuf_size2_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_27_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_28_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_29_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_136_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_30_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_31_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_143_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_32_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_33_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_159 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_150_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_34_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_35_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_157_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_36_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_179 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_37_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_195 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_164_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_38_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_197 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_39_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_18__0_ -----

//----- Default net type -----
`default_nettype wire



