//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Connection Blocks[6][5]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jul  5 01:26:08 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for cbx_6__5_ -----
module cbx_6__5_(prog_clk,
                 chanx_left_in,
                 chanx_right_in,
                 ccff_head,
                 chanx_left_out,
                 chanx_right_out,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_reset_0_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_0_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_1_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_2_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_3_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_4_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_5_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_6_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_7_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_8_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_9_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_10_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_11_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_12_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_13_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_14_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_15_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_16_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_17_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_18_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_19_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_20_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_21_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_22_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_23_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_24_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_25_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_26_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_27_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_28_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_29_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_30_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_31_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_32_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_33_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_34_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_35_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_36_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_37_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_38_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_39_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_40_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_41_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_42_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_43_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_44_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_45_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_46_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_47_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_48_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_49_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_50_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_51_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_52_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_53_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_54_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_55_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_56_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_57_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_58_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_59_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_60_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_61_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_62_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_63_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_64_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_65_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_66_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_67_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_68_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_69_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_0_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_1_,
                 top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_2_,
                 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_,
                 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_,
                 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:284] chanx_left_in;
//----- INPUT PORTS -----
input [0:284] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:284] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:284] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_0_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_1_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_2_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_3_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_4_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_5_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_6_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_7_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_8_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_9_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_10_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_11_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_12_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_13_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_14_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_15_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_16_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_17_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_18_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_19_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_20_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_21_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_22_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_23_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_24_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_25_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_26_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_27_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_28_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_29_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_30_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_31_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_32_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_33_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_34_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_35_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_36_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_37_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_38_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_39_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_40_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_41_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_42_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_43_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_44_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_45_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_46_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_47_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_48_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_49_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_50_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_51_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_52_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_53_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_54_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_55_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_56_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_57_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_58_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_59_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_60_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_61_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_62_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_63_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_64_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_65_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_66_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_67_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_68_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_69_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_0_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_1_;
//----- OUTPUT PORTS -----
output [0:0] top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:6] mux_tree_tapbuf_size96_0_sram;
wire [0:6] mux_tree_tapbuf_size96_0_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_10_sram;
wire [0:6] mux_tree_tapbuf_size96_10_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_11_sram;
wire [0:6] mux_tree_tapbuf_size96_11_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_12_sram;
wire [0:6] mux_tree_tapbuf_size96_12_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_13_sram;
wire [0:6] mux_tree_tapbuf_size96_13_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_14_sram;
wire [0:6] mux_tree_tapbuf_size96_14_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_15_sram;
wire [0:6] mux_tree_tapbuf_size96_15_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_16_sram;
wire [0:6] mux_tree_tapbuf_size96_16_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_17_sram;
wire [0:6] mux_tree_tapbuf_size96_17_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_18_sram;
wire [0:6] mux_tree_tapbuf_size96_18_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_19_sram;
wire [0:6] mux_tree_tapbuf_size96_19_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_1_sram;
wire [0:6] mux_tree_tapbuf_size96_1_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_20_sram;
wire [0:6] mux_tree_tapbuf_size96_20_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_21_sram;
wire [0:6] mux_tree_tapbuf_size96_21_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_22_sram;
wire [0:6] mux_tree_tapbuf_size96_22_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_23_sram;
wire [0:6] mux_tree_tapbuf_size96_23_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_24_sram;
wire [0:6] mux_tree_tapbuf_size96_24_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_25_sram;
wire [0:6] mux_tree_tapbuf_size96_25_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_26_sram;
wire [0:6] mux_tree_tapbuf_size96_26_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_27_sram;
wire [0:6] mux_tree_tapbuf_size96_27_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_28_sram;
wire [0:6] mux_tree_tapbuf_size96_28_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_29_sram;
wire [0:6] mux_tree_tapbuf_size96_29_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_2_sram;
wire [0:6] mux_tree_tapbuf_size96_2_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_30_sram;
wire [0:6] mux_tree_tapbuf_size96_30_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_31_sram;
wire [0:6] mux_tree_tapbuf_size96_31_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_32_sram;
wire [0:6] mux_tree_tapbuf_size96_32_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_33_sram;
wire [0:6] mux_tree_tapbuf_size96_33_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_34_sram;
wire [0:6] mux_tree_tapbuf_size96_34_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_35_sram;
wire [0:6] mux_tree_tapbuf_size96_35_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_36_sram;
wire [0:6] mux_tree_tapbuf_size96_36_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_37_sram;
wire [0:6] mux_tree_tapbuf_size96_37_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_38_sram;
wire [0:6] mux_tree_tapbuf_size96_38_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_39_sram;
wire [0:6] mux_tree_tapbuf_size96_39_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_3_sram;
wire [0:6] mux_tree_tapbuf_size96_3_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_40_sram;
wire [0:6] mux_tree_tapbuf_size96_40_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_41_sram;
wire [0:6] mux_tree_tapbuf_size96_41_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_42_sram;
wire [0:6] mux_tree_tapbuf_size96_42_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_43_sram;
wire [0:6] mux_tree_tapbuf_size96_43_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_44_sram;
wire [0:6] mux_tree_tapbuf_size96_44_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_45_sram;
wire [0:6] mux_tree_tapbuf_size96_45_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_46_sram;
wire [0:6] mux_tree_tapbuf_size96_46_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_47_sram;
wire [0:6] mux_tree_tapbuf_size96_47_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_48_sram;
wire [0:6] mux_tree_tapbuf_size96_48_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_49_sram;
wire [0:6] mux_tree_tapbuf_size96_49_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_4_sram;
wire [0:6] mux_tree_tapbuf_size96_4_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_50_sram;
wire [0:6] mux_tree_tapbuf_size96_50_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_51_sram;
wire [0:6] mux_tree_tapbuf_size96_51_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_52_sram;
wire [0:6] mux_tree_tapbuf_size96_52_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_53_sram;
wire [0:6] mux_tree_tapbuf_size96_53_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_54_sram;
wire [0:6] mux_tree_tapbuf_size96_54_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_55_sram;
wire [0:6] mux_tree_tapbuf_size96_55_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_56_sram;
wire [0:6] mux_tree_tapbuf_size96_56_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_57_sram;
wire [0:6] mux_tree_tapbuf_size96_57_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_58_sram;
wire [0:6] mux_tree_tapbuf_size96_58_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_59_sram;
wire [0:6] mux_tree_tapbuf_size96_59_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_5_sram;
wire [0:6] mux_tree_tapbuf_size96_5_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_60_sram;
wire [0:6] mux_tree_tapbuf_size96_60_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_61_sram;
wire [0:6] mux_tree_tapbuf_size96_61_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_62_sram;
wire [0:6] mux_tree_tapbuf_size96_62_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_63_sram;
wire [0:6] mux_tree_tapbuf_size96_63_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_64_sram;
wire [0:6] mux_tree_tapbuf_size96_64_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_65_sram;
wire [0:6] mux_tree_tapbuf_size96_65_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_66_sram;
wire [0:6] mux_tree_tapbuf_size96_66_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_67_sram;
wire [0:6] mux_tree_tapbuf_size96_67_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_68_sram;
wire [0:6] mux_tree_tapbuf_size96_68_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_69_sram;
wire [0:6] mux_tree_tapbuf_size96_69_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_6_sram;
wire [0:6] mux_tree_tapbuf_size96_6_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_70_sram;
wire [0:6] mux_tree_tapbuf_size96_70_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_71_sram;
wire [0:6] mux_tree_tapbuf_size96_71_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_72_sram;
wire [0:6] mux_tree_tapbuf_size96_72_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_73_sram;
wire [0:6] mux_tree_tapbuf_size96_73_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_74_sram;
wire [0:6] mux_tree_tapbuf_size96_74_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_75_sram;
wire [0:6] mux_tree_tapbuf_size96_75_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_76_sram;
wire [0:6] mux_tree_tapbuf_size96_76_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_7_sram;
wire [0:6] mux_tree_tapbuf_size96_7_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_8_sram;
wire [0:6] mux_tree_tapbuf_size96_8_sram_inv;
wire [0:6] mux_tree_tapbuf_size96_9_sram;
wire [0:6] mux_tree_tapbuf_size96_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size96_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size96_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[0] = chanx_left_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[1] = chanx_left_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[2] = chanx_left_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[3] = chanx_left_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[4] = chanx_left_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[5] = chanx_left_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[6] = chanx_left_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[7] = chanx_left_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[8] = chanx_left_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[9] = chanx_left_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[10] = chanx_left_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[11] = chanx_left_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[12] = chanx_left_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[13] = chanx_left_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[14] = chanx_left_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[15] = chanx_left_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[16] = chanx_left_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chanx_left_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[18] = chanx_left_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[19] = chanx_left_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[20] = chanx_left_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[21] = chanx_left_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[22] = chanx_left_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[23] = chanx_left_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[24] = chanx_left_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[25] = chanx_left_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[26] = chanx_left_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[27] = chanx_left_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[28] = chanx_left_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[29] = chanx_left_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[30] = chanx_left_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[31] = chanx_left_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[32] = chanx_left_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[33] = chanx_left_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[34] = chanx_left_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[35] = chanx_left_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[36] = chanx_left_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[37] = chanx_left_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[38] = chanx_left_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[39] = chanx_left_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[40] = chanx_left_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[41] = chanx_left_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[42] = chanx_left_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[43] = chanx_left_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[44] = chanx_left_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[45] = chanx_left_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[46] = chanx_left_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[47] = chanx_left_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[48] = chanx_left_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[49] = chanx_left_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[50] = chanx_left_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[51] = chanx_left_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[52] = chanx_left_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[53] = chanx_left_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[54] = chanx_left_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[55] = chanx_left_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[56] = chanx_left_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[57] = chanx_left_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[58] = chanx_left_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[59] = chanx_left_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[60] = chanx_left_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[61] = chanx_left_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[62] = chanx_left_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[63] = chanx_left_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[64] = chanx_left_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[65] = chanx_left_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[66] = chanx_left_in[66];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[67] = chanx_left_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[68] = chanx_left_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[69] = chanx_left_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[70] = chanx_left_in[70];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[71] = chanx_left_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[72] = chanx_left_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[73] = chanx_left_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[74] = chanx_left_in[74];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[75] = chanx_left_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[76] = chanx_left_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[77] = chanx_left_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[78] = chanx_left_in[78];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[79] = chanx_left_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[80] = chanx_left_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[81] = chanx_left_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[82] = chanx_left_in[82];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[83] = chanx_left_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[84] = chanx_left_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[85] = chanx_left_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[86] = chanx_left_in[86];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[87] = chanx_left_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[88] = chanx_left_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[89] = chanx_left_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[90] = chanx_left_in[90];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[91] = chanx_left_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[92] = chanx_left_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[93] = chanx_left_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[94] = chanx_left_in[94];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[95] = chanx_left_in[95];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[96] = chanx_left_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[97] = chanx_left_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[98] = chanx_left_in[98];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[99] = chanx_left_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[100] = chanx_left_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[101] = chanx_left_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[102] = chanx_left_in[102];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[103] = chanx_left_in[103];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[104] = chanx_left_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[105] = chanx_left_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[106] = chanx_left_in[106];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[107] = chanx_left_in[107];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[108] = chanx_left_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[109] = chanx_left_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[110] = chanx_left_in[110];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[111] = chanx_left_in[111];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[112] = chanx_left_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[113] = chanx_left_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[114] = chanx_left_in[114];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[115] = chanx_left_in[115];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[116] = chanx_left_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[117] = chanx_left_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[118] = chanx_left_in[118];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[119] = chanx_left_in[119];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[120] = chanx_left_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[121] = chanx_left_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[122] = chanx_left_in[122];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[123] = chanx_left_in[123];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[124] = chanx_left_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[125] = chanx_left_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[126] = chanx_left_in[126];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[127] = chanx_left_in[127];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[128] = chanx_left_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[129] = chanx_left_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[130] = chanx_left_in[130];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[131] = chanx_left_in[131];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[132] = chanx_left_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[133] = chanx_left_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[134] = chanx_left_in[134];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[135] = chanx_left_in[135];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[136] = chanx_left_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[137] = chanx_left_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[138] = chanx_left_in[138];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[139] = chanx_left_in[139];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[140] = chanx_left_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[141] = chanx_left_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[142] = chanx_left_in[142];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[143] = chanx_left_in[143];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[144] = chanx_left_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[145] = chanx_left_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[146] = chanx_left_in[146];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[147] = chanx_left_in[147];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[148] = chanx_left_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[149] = chanx_left_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[150] = chanx_left_in[150];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[151] = chanx_left_in[151];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[152] = chanx_left_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[153] = chanx_left_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[154] = chanx_left_in[154];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[155] = chanx_left_in[155];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[156] = chanx_left_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[157] = chanx_left_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[158] = chanx_left_in[158];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[159] = chanx_left_in[159];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[160] = chanx_left_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[161] = chanx_left_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[162] = chanx_left_in[162];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[163] = chanx_left_in[163];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[164] = chanx_left_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[165] = chanx_left_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[166] = chanx_left_in[166];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[167] = chanx_left_in[167];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[168] = chanx_left_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[169] = chanx_left_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[170] = chanx_left_in[170];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[171] = chanx_left_in[171];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[172] = chanx_left_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[173] = chanx_left_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[174] = chanx_left_in[174];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[175] = chanx_left_in[175];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[176] = chanx_left_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[177] = chanx_left_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[178] = chanx_left_in[178];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[179] = chanx_left_in[179];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[180] = chanx_left_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[181] = chanx_left_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[182] = chanx_left_in[182];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[183] = chanx_left_in[183];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[184] = chanx_left_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[185] = chanx_left_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[186] = chanx_left_in[186];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[187] = chanx_left_in[187];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[188] = chanx_left_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[189] = chanx_left_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[190] = chanx_left_in[190];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[191] = chanx_left_in[191];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[192] = chanx_left_in[192];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[193] = chanx_left_in[193];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[194] = chanx_left_in[194];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[195] = chanx_left_in[195];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[196] = chanx_left_in[196];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[197] = chanx_left_in[197];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[198] = chanx_left_in[198];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[199] = chanx_left_in[199];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[200] = chanx_left_in[200];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[201] = chanx_left_in[201];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[202] = chanx_left_in[202];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[203] = chanx_left_in[203];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[204] = chanx_left_in[204];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[205] = chanx_left_in[205];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[206] = chanx_left_in[206];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[207] = chanx_left_in[207];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[208] = chanx_left_in[208];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[209] = chanx_left_in[209];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[210] = chanx_left_in[210];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[211] = chanx_left_in[211];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[212] = chanx_left_in[212];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[213] = chanx_left_in[213];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[214] = chanx_left_in[214];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[215] = chanx_left_in[215];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[216] = chanx_left_in[216];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[217] = chanx_left_in[217];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[218] = chanx_left_in[218];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[219] = chanx_left_in[219];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[220] = chanx_left_in[220];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[221] = chanx_left_in[221];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[222] = chanx_left_in[222];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[223] = chanx_left_in[223];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[224] = chanx_left_in[224];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[225] = chanx_left_in[225];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[226] = chanx_left_in[226];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[227] = chanx_left_in[227];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[228] = chanx_left_in[228];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[229] = chanx_left_in[229];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[230] = chanx_left_in[230];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[231] = chanx_left_in[231];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[232] = chanx_left_in[232];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[233] = chanx_left_in[233];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[234] = chanx_left_in[234];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[235] = chanx_left_in[235];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[236] = chanx_left_in[236];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[237] = chanx_left_in[237];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[238] = chanx_left_in[238];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[239] = chanx_left_in[239];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[240] = chanx_left_in[240];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[241] = chanx_left_in[241];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[242] = chanx_left_in[242];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[243] = chanx_left_in[243];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[244] = chanx_left_in[244];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[245] = chanx_left_in[245];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[246] = chanx_left_in[246];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[247] = chanx_left_in[247];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[248] = chanx_left_in[248];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[249] = chanx_left_in[249];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[250] = chanx_left_in[250];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[251] = chanx_left_in[251];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[252] = chanx_left_in[252];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[253] = chanx_left_in[253];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[254] = chanx_left_in[254];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[255] = chanx_left_in[255];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[256] = chanx_left_in[256];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[257] = chanx_left_in[257];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[258] = chanx_left_in[258];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[259] = chanx_left_in[259];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[260] = chanx_left_in[260];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[261] = chanx_left_in[261];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[262] = chanx_left_in[262];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[263] = chanx_left_in[263];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[264] = chanx_left_in[264];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[265] = chanx_left_in[265];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[266] = chanx_left_in[266];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[267] = chanx_left_in[267];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[268] = chanx_left_in[268];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[269] = chanx_left_in[269];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[270] = chanx_left_in[270];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[271] = chanx_left_in[271];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[272] = chanx_left_in[272];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[273] = chanx_left_in[273];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[274] = chanx_left_in[274];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[275] = chanx_left_in[275];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[276] = chanx_left_in[276];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[277] = chanx_left_in[277];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[278] = chanx_left_in[278];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[279] = chanx_left_in[279];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[280] = chanx_left_in[280];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[281] = chanx_left_in[281];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[282] = chanx_left_in[282];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[283] = chanx_left_in[283];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[284] = chanx_left_in[284];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[0] = chanx_right_in[0];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[1] = chanx_right_in[1];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[2] = chanx_right_in[2];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[3] = chanx_right_in[3];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[4] = chanx_right_in[4];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[5] = chanx_right_in[5];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[6] = chanx_right_in[6];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[7] = chanx_right_in[7];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[8] = chanx_right_in[8];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[9] = chanx_right_in[9];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[10] = chanx_right_in[10];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[11] = chanx_right_in[11];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[12] = chanx_right_in[12];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[13] = chanx_right_in[13];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[14] = chanx_right_in[14];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[15] = chanx_right_in[15];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[16] = chanx_right_in[16];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[17] = chanx_right_in[17];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[18] = chanx_right_in[18];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[19] = chanx_right_in[19];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[20] = chanx_right_in[20];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[21] = chanx_right_in[21];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[22] = chanx_right_in[22];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[23] = chanx_right_in[23];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[24] = chanx_right_in[24];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[25] = chanx_right_in[25];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[26] = chanx_right_in[26];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[27] = chanx_right_in[27];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[28] = chanx_right_in[28];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[29] = chanx_right_in[29];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[30] = chanx_right_in[30];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[31] = chanx_right_in[31];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[32] = chanx_right_in[32];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[33] = chanx_right_in[33];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[34] = chanx_right_in[34];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[35] = chanx_right_in[35];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[36] = chanx_right_in[36];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[37] = chanx_right_in[37];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[38] = chanx_right_in[38];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[39] = chanx_right_in[39];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[40] = chanx_right_in[40];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[41] = chanx_right_in[41];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[42] = chanx_right_in[42];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[43] = chanx_right_in[43];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[44] = chanx_right_in[44];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[45] = chanx_right_in[45];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[46] = chanx_right_in[46];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[47] = chanx_right_in[47];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[48] = chanx_right_in[48];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[49] = chanx_right_in[49];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[50] = chanx_right_in[50];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[51] = chanx_right_in[51];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[52] = chanx_right_in[52];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[53] = chanx_right_in[53];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[54] = chanx_right_in[54];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[55] = chanx_right_in[55];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[56] = chanx_right_in[56];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[57] = chanx_right_in[57];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[58] = chanx_right_in[58];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[59] = chanx_right_in[59];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[60] = chanx_right_in[60];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[61] = chanx_right_in[61];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[62] = chanx_right_in[62];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[63] = chanx_right_in[63];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[64] = chanx_right_in[64];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[65] = chanx_right_in[65];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[66] = chanx_right_in[66];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[67] = chanx_right_in[67];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[68] = chanx_right_in[68];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[69] = chanx_right_in[69];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[70] = chanx_right_in[70];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[71] = chanx_right_in[71];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[72] = chanx_right_in[72];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[73] = chanx_right_in[73];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[74] = chanx_right_in[74];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[75] = chanx_right_in[75];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[76] = chanx_right_in[76];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[77] = chanx_right_in[77];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[78] = chanx_right_in[78];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[79] = chanx_right_in[79];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[80] = chanx_right_in[80];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[81] = chanx_right_in[81];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[82] = chanx_right_in[82];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[83] = chanx_right_in[83];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[84] = chanx_right_in[84];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[85] = chanx_right_in[85];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[86] = chanx_right_in[86];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[87] = chanx_right_in[87];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[88] = chanx_right_in[88];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[89] = chanx_right_in[89];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[90] = chanx_right_in[90];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[91] = chanx_right_in[91];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[92] = chanx_right_in[92];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[93] = chanx_right_in[93];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[94] = chanx_right_in[94];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[95] = chanx_right_in[95];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[96] = chanx_right_in[96];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[97] = chanx_right_in[97];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[98] = chanx_right_in[98];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[99] = chanx_right_in[99];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[100] = chanx_right_in[100];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[101] = chanx_right_in[101];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[102] = chanx_right_in[102];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[103] = chanx_right_in[103];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[104] = chanx_right_in[104];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[105] = chanx_right_in[105];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[106] = chanx_right_in[106];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[107] = chanx_right_in[107];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[108] = chanx_right_in[108];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[109] = chanx_right_in[109];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[110] = chanx_right_in[110];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[111] = chanx_right_in[111];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[112] = chanx_right_in[112];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[113] = chanx_right_in[113];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[114] = chanx_right_in[114];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[115] = chanx_right_in[115];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[116] = chanx_right_in[116];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[117] = chanx_right_in[117];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[118] = chanx_right_in[118];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[119] = chanx_right_in[119];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[120] = chanx_right_in[120];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[121] = chanx_right_in[121];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[122] = chanx_right_in[122];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[123] = chanx_right_in[123];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[124] = chanx_right_in[124];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[125] = chanx_right_in[125];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[126] = chanx_right_in[126];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[127] = chanx_right_in[127];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[128] = chanx_right_in[128];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[129] = chanx_right_in[129];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[130] = chanx_right_in[130];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[131] = chanx_right_in[131];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[132] = chanx_right_in[132];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[133] = chanx_right_in[133];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[134] = chanx_right_in[134];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[135] = chanx_right_in[135];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[136] = chanx_right_in[136];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[137] = chanx_right_in[137];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[138] = chanx_right_in[138];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[139] = chanx_right_in[139];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[140] = chanx_right_in[140];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[141] = chanx_right_in[141];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[142] = chanx_right_in[142];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[143] = chanx_right_in[143];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[144] = chanx_right_in[144];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[145] = chanx_right_in[145];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[146] = chanx_right_in[146];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[147] = chanx_right_in[147];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[148] = chanx_right_in[148];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[149] = chanx_right_in[149];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[150] = chanx_right_in[150];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[151] = chanx_right_in[151];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[152] = chanx_right_in[152];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[153] = chanx_right_in[153];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[154] = chanx_right_in[154];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[155] = chanx_right_in[155];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[156] = chanx_right_in[156];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[157] = chanx_right_in[157];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[158] = chanx_right_in[158];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[159] = chanx_right_in[159];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[160] = chanx_right_in[160];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[161] = chanx_right_in[161];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[162] = chanx_right_in[162];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[163] = chanx_right_in[163];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[164] = chanx_right_in[164];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[165] = chanx_right_in[165];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[166] = chanx_right_in[166];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[167] = chanx_right_in[167];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[168] = chanx_right_in[168];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[169] = chanx_right_in[169];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[170] = chanx_right_in[170];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[171] = chanx_right_in[171];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[172] = chanx_right_in[172];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[173] = chanx_right_in[173];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[174] = chanx_right_in[174];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[175] = chanx_right_in[175];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[176] = chanx_right_in[176];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[177] = chanx_right_in[177];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[178] = chanx_right_in[178];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[179] = chanx_right_in[179];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[180] = chanx_right_in[180];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[181] = chanx_right_in[181];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[182] = chanx_right_in[182];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[183] = chanx_right_in[183];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[184] = chanx_right_in[184];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[185] = chanx_right_in[185];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[186] = chanx_right_in[186];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[187] = chanx_right_in[187];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[188] = chanx_right_in[188];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[189] = chanx_right_in[189];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[190] = chanx_right_in[190];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[191] = chanx_right_in[191];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[192] = chanx_right_in[192];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[193] = chanx_right_in[193];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[194] = chanx_right_in[194];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[195] = chanx_right_in[195];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[196] = chanx_right_in[196];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[197] = chanx_right_in[197];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[198] = chanx_right_in[198];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[199] = chanx_right_in[199];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[200] = chanx_right_in[200];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[201] = chanx_right_in[201];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[202] = chanx_right_in[202];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[203] = chanx_right_in[203];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[204] = chanx_right_in[204];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[205] = chanx_right_in[205];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[206] = chanx_right_in[206];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[207] = chanx_right_in[207];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[208] = chanx_right_in[208];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[209] = chanx_right_in[209];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[210] = chanx_right_in[210];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[211] = chanx_right_in[211];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[212] = chanx_right_in[212];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[213] = chanx_right_in[213];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[214] = chanx_right_in[214];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[215] = chanx_right_in[215];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[216] = chanx_right_in[216];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[217] = chanx_right_in[217];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[218] = chanx_right_in[218];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[219] = chanx_right_in[219];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[220] = chanx_right_in[220];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[221] = chanx_right_in[221];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[222] = chanx_right_in[222];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[223] = chanx_right_in[223];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[224] = chanx_right_in[224];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[225] = chanx_right_in[225];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[226] = chanx_right_in[226];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[227] = chanx_right_in[227];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[228] = chanx_right_in[228];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[229] = chanx_right_in[229];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[230] = chanx_right_in[230];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[231] = chanx_right_in[231];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[232] = chanx_right_in[232];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[233] = chanx_right_in[233];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[234] = chanx_right_in[234];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[235] = chanx_right_in[235];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[236] = chanx_right_in[236];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[237] = chanx_right_in[237];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[238] = chanx_right_in[238];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[239] = chanx_right_in[239];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[240] = chanx_right_in[240];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[241] = chanx_right_in[241];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[242] = chanx_right_in[242];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[243] = chanx_right_in[243];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[244] = chanx_right_in[244];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[245] = chanx_right_in[245];
// ----- Local connection due to Wire 531 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[246] = chanx_right_in[246];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[247] = chanx_right_in[247];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[248] = chanx_right_in[248];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[249] = chanx_right_in[249];
// ----- Local connection due to Wire 535 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[250] = chanx_right_in[250];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[251] = chanx_right_in[251];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[252] = chanx_right_in[252];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[253] = chanx_right_in[253];
// ----- Local connection due to Wire 539 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[254] = chanx_right_in[254];
// ----- Local connection due to Wire 540 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[255] = chanx_right_in[255];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[256] = chanx_right_in[256];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[257] = chanx_right_in[257];
// ----- Local connection due to Wire 543 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[258] = chanx_right_in[258];
// ----- Local connection due to Wire 544 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[259] = chanx_right_in[259];
// ----- Local connection due to Wire 545 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[260] = chanx_right_in[260];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[261] = chanx_right_in[261];
// ----- Local connection due to Wire 547 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[262] = chanx_right_in[262];
// ----- Local connection due to Wire 548 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[263] = chanx_right_in[263];
// ----- Local connection due to Wire 549 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[264] = chanx_right_in[264];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[265] = chanx_right_in[265];
// ----- Local connection due to Wire 551 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[266] = chanx_right_in[266];
// ----- Local connection due to Wire 552 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[267] = chanx_right_in[267];
// ----- Local connection due to Wire 553 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[268] = chanx_right_in[268];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[269] = chanx_right_in[269];
// ----- Local connection due to Wire 555 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[270] = chanx_right_in[270];
// ----- Local connection due to Wire 556 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[271] = chanx_right_in[271];
// ----- Local connection due to Wire 557 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[272] = chanx_right_in[272];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[273] = chanx_right_in[273];
// ----- Local connection due to Wire 559 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[274] = chanx_right_in[274];
// ----- Local connection due to Wire 560 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[275] = chanx_right_in[275];
// ----- Local connection due to Wire 561 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[276] = chanx_right_in[276];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[277] = chanx_right_in[277];
// ----- Local connection due to Wire 563 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[278] = chanx_right_in[278];
// ----- Local connection due to Wire 564 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[279] = chanx_right_in[279];
// ----- Local connection due to Wire 565 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[280] = chanx_right_in[280];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[281] = chanx_right_in[281];
// ----- Local connection due to Wire 567 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[282] = chanx_right_in[282];
// ----- Local connection due to Wire 568 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[283] = chanx_right_in[283];
// ----- Local connection due to Wire 569 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[284] = chanx_right_in[284];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size96 mux_bottom_ipin_0 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_0_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_0_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_reset_0_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_1 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_1_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_1_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_0_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_2 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_2_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_2_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_1_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_3 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_3_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_3_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_2_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_4 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_4_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_4_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_3_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_5 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_5_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_5_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_4_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_6 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_6_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_6_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_5_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_7 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_7_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_7_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_6_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_8 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_8_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_8_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_7_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_9 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_9_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_9_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_8_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_10 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_10_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_10_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_9_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_11 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_11_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_11_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_10_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_12 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_12_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_12_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_11_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_13 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_13_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_13_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_12_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_14 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_14_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_14_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_13_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_15 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_15_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_15_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_14_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_16 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_16_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_16_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_15_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_17 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_17_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_17_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_16_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_18 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_18_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_18_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_17_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_19 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_19_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_19_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_18_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_20 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_20_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_20_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_19_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_21 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_21_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_21_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_20_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_22 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_22_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_22_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_21_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_23 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_23_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_23_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_22_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_24 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_24_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_24_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_23_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_25 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_25_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_25_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_24_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_26 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_26_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_26_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_25_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_27 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_27_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_27_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_26_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_28 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_28_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_28_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_27_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_29 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_29_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_29_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_28_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_30 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_30_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_30_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_29_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_31 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_31_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_31_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_30_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_32 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_32_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_32_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_31_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_33 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_33_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_33_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_32_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_34 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_34_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_34_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_33_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_35 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_35_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_35_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_34_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_36 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_36_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_36_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_35_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_37 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_37_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_37_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_36_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_38 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_38_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_38_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_37_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_39 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_39_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_39_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_38_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_40 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_40_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_40_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_39_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_41 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_41_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_41_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_40_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_42 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_42_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_42_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_41_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_43 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_43_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_43_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_42_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_44 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_44_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_44_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_43_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_45 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_45_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_45_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_44_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_46 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_46_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_46_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_45_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_47 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_47_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_47_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_46_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_48 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_48_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_48_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_47_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_49 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_49_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_49_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_48_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_50 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_50_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_50_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_49_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_51 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_51_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_51_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_50_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_52 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_52_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_52_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_51_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_53 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_53_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_53_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_52_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_54 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_54_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_54_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_53_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_55 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_55_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_55_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_54_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_56 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_56_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_56_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_55_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_57 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_57_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_57_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_56_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_58 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_58_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_58_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_57_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_59 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_59_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_59_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_58_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_60 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_60_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_60_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_59_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_61 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_61_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_61_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_60_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_62 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_62_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_62_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_61_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_63 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_63_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_63_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_62_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_64 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_64_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_64_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_63_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_65 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_65_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_65_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_64_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_66 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_66_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_66_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_65_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_67 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_67_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_67_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_66_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_68 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[68], chanx_right_in[68], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_68_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_68_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_67_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_69 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[69], chanx_right_in[69], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_69_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_69_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_68_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_70 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[70], chanx_right_in[70], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_70_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_70_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_2_69_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_71 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[8], chanx_right_in[8], chanx_left_in[14], chanx_right_in[14], chanx_left_in[20], chanx_right_in[20], chanx_left_in[26], chanx_right_in[26], chanx_left_in[32], chanx_right_in[32], chanx_left_in[38], chanx_right_in[38], chanx_left_in[44], chanx_right_in[44], chanx_left_in[50], chanx_right_in[50], chanx_left_in[56], chanx_right_in[56], chanx_left_in[62], chanx_right_in[62], chanx_left_in[68], chanx_right_in[68], chanx_left_in[71], chanx_right_in[71], chanx_left_in[77], chanx_right_in[77], chanx_left_in[83], chanx_right_in[83], chanx_left_in[89], chanx_right_in[89], chanx_left_in[95], chanx_right_in[95], chanx_left_in[101], chanx_right_in[101], chanx_left_in[107], chanx_right_in[107], chanx_left_in[113], chanx_right_in[113], chanx_left_in[119], chanx_right_in[119], chanx_left_in[125], chanx_right_in[125], chanx_left_in[131], chanx_right_in[131], chanx_left_in[137], chanx_right_in[137], chanx_left_in[143], chanx_right_in[143], chanx_left_in[149], chanx_right_in[149], chanx_left_in[155], chanx_right_in[155], chanx_left_in[161], chanx_right_in[161], chanx_left_in[167], chanx_right_in[167], chanx_left_in[173], chanx_right_in[173], chanx_left_in[179], chanx_right_in[179], chanx_left_in[185], chanx_right_in[185], chanx_left_in[191], chanx_right_in[191], chanx_left_in[197], chanx_right_in[197], chanx_left_in[203], chanx_right_in[203], chanx_left_in[209], chanx_right_in[209], chanx_left_in[215], chanx_right_in[215], chanx_left_in[221], chanx_right_in[221], chanx_left_in[227], chanx_right_in[227], chanx_left_in[233], chanx_right_in[233], chanx_left_in[239], chanx_right_in[239], chanx_left_in[245], chanx_right_in[245], chanx_left_in[251], chanx_right_in[251], chanx_left_in[257], chanx_right_in[257], chanx_left_in[263], chanx_right_in[263], chanx_left_in[269], chanx_right_in[269], chanx_left_in[275], chanx_right_in[275], chanx_left_in[281], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size96_71_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_71_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_0_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_72 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[9], chanx_right_in[9], chanx_left_in[15], chanx_right_in[15], chanx_left_in[21], chanx_right_in[21], chanx_left_in[27], chanx_right_in[27], chanx_left_in[33], chanx_right_in[33], chanx_left_in[39], chanx_right_in[39], chanx_left_in[45], chanx_right_in[45], chanx_left_in[51], chanx_right_in[51], chanx_left_in[57], chanx_right_in[57], chanx_left_in[63], chanx_right_in[63], chanx_left_in[69], chanx_right_in[69], chanx_left_in[72], chanx_right_in[72], chanx_left_in[78], chanx_right_in[78], chanx_left_in[84], chanx_right_in[84], chanx_left_in[90], chanx_right_in[90], chanx_left_in[96], chanx_right_in[96], chanx_left_in[102], chanx_right_in[102], chanx_left_in[108], chanx_right_in[108], chanx_left_in[114], chanx_right_in[114], chanx_left_in[120], chanx_right_in[120], chanx_left_in[126], chanx_right_in[126], chanx_left_in[132], chanx_right_in[132], chanx_left_in[138], chanx_right_in[138], chanx_left_in[144], chanx_right_in[144], chanx_left_in[150], chanx_right_in[150], chanx_left_in[156], chanx_right_in[156], chanx_left_in[162], chanx_right_in[162], chanx_left_in[168], chanx_right_in[168], chanx_left_in[174], chanx_right_in[174], chanx_left_in[180], chanx_right_in[180], chanx_left_in[186], chanx_right_in[186], chanx_left_in[192], chanx_right_in[192], chanx_left_in[198], chanx_right_in[198], chanx_left_in[204], chanx_right_in[204], chanx_left_in[210], chanx_right_in[210], chanx_left_in[216], chanx_right_in[216], chanx_left_in[222], chanx_right_in[222], chanx_left_in[228], chanx_right_in[228], chanx_left_in[234], chanx_right_in[234], chanx_left_in[240], chanx_right_in[240], chanx_left_in[246], chanx_right_in[246], chanx_left_in[252], chanx_right_in[252], chanx_left_in[258], chanx_right_in[258], chanx_left_in[264], chanx_right_in[264], chanx_left_in[270], chanx_right_in[270], chanx_left_in[276], chanx_right_in[276], chanx_left_in[282], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size96_72_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_72_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_1_));

	mux_tree_tapbuf_size96 mux_bottom_ipin_73 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[10], chanx_right_in[10], chanx_left_in[16], chanx_right_in[16], chanx_left_in[22], chanx_right_in[22], chanx_left_in[28], chanx_right_in[28], chanx_left_in[34], chanx_right_in[34], chanx_left_in[40], chanx_right_in[40], chanx_left_in[46], chanx_right_in[46], chanx_left_in[52], chanx_right_in[52], chanx_left_in[58], chanx_right_in[58], chanx_left_in[64], chanx_right_in[64], chanx_left_in[70], chanx_right_in[70], chanx_left_in[73], chanx_right_in[73], chanx_left_in[79], chanx_right_in[79], chanx_left_in[85], chanx_right_in[85], chanx_left_in[91], chanx_right_in[91], chanx_left_in[97], chanx_right_in[97], chanx_left_in[103], chanx_right_in[103], chanx_left_in[109], chanx_right_in[109], chanx_left_in[115], chanx_right_in[115], chanx_left_in[121], chanx_right_in[121], chanx_left_in[127], chanx_right_in[127], chanx_left_in[133], chanx_right_in[133], chanx_left_in[139], chanx_right_in[139], chanx_left_in[145], chanx_right_in[145], chanx_left_in[151], chanx_right_in[151], chanx_left_in[157], chanx_right_in[157], chanx_left_in[163], chanx_right_in[163], chanx_left_in[169], chanx_right_in[169], chanx_left_in[175], chanx_right_in[175], chanx_left_in[181], chanx_right_in[181], chanx_left_in[187], chanx_right_in[187], chanx_left_in[193], chanx_right_in[193], chanx_left_in[199], chanx_right_in[199], chanx_left_in[205], chanx_right_in[205], chanx_left_in[211], chanx_right_in[211], chanx_left_in[217], chanx_right_in[217], chanx_left_in[223], chanx_right_in[223], chanx_left_in[229], chanx_right_in[229], chanx_left_in[235], chanx_right_in[235], chanx_left_in[241], chanx_right_in[241], chanx_left_in[247], chanx_right_in[247], chanx_left_in[253], chanx_right_in[253], chanx_left_in[259], chanx_right_in[259], chanx_left_in[265], chanx_right_in[265], chanx_left_in[271], chanx_right_in[271], chanx_left_in[277], chanx_right_in[277], chanx_left_in[283], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size96_73_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_73_sram_inv[0:6]),
		.out(top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_2_));

	mux_tree_tapbuf_size96 mux_top_ipin_0 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[11], chanx_right_in[11], chanx_left_in[17], chanx_right_in[17], chanx_left_in[23], chanx_right_in[23], chanx_left_in[29], chanx_right_in[29], chanx_left_in[35], chanx_right_in[35], chanx_left_in[41], chanx_right_in[41], chanx_left_in[47], chanx_right_in[47], chanx_left_in[53], chanx_right_in[53], chanx_left_in[59], chanx_right_in[59], chanx_left_in[65], chanx_right_in[65], chanx_left_in[71], chanx_right_in[71], chanx_left_in[74], chanx_right_in[74], chanx_left_in[80], chanx_right_in[80], chanx_left_in[86], chanx_right_in[86], chanx_left_in[92], chanx_right_in[92], chanx_left_in[98], chanx_right_in[98], chanx_left_in[104], chanx_right_in[104], chanx_left_in[110], chanx_right_in[110], chanx_left_in[116], chanx_right_in[116], chanx_left_in[122], chanx_right_in[122], chanx_left_in[128], chanx_right_in[128], chanx_left_in[134], chanx_right_in[134], chanx_left_in[140], chanx_right_in[140], chanx_left_in[146], chanx_right_in[146], chanx_left_in[152], chanx_right_in[152], chanx_left_in[158], chanx_right_in[158], chanx_left_in[164], chanx_right_in[164], chanx_left_in[170], chanx_right_in[170], chanx_left_in[176], chanx_right_in[176], chanx_left_in[182], chanx_right_in[182], chanx_left_in[188], chanx_right_in[188], chanx_left_in[194], chanx_right_in[194], chanx_left_in[200], chanx_right_in[200], chanx_left_in[206], chanx_right_in[206], chanx_left_in[212], chanx_right_in[212], chanx_left_in[218], chanx_right_in[218], chanx_left_in[224], chanx_right_in[224], chanx_left_in[230], chanx_right_in[230], chanx_left_in[236], chanx_right_in[236], chanx_left_in[242], chanx_right_in[242], chanx_left_in[248], chanx_right_in[248], chanx_left_in[254], chanx_right_in[254], chanx_left_in[260], chanx_right_in[260], chanx_left_in[266], chanx_right_in[266], chanx_left_in[272], chanx_right_in[272], chanx_left_in[278], chanx_right_in[278], chanx_left_in[284], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size96_74_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_74_sram_inv[0:6]),
		.out(bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_));

	mux_tree_tapbuf_size96 mux_top_ipin_1 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[6], chanx_right_in[6], chanx_left_in[12], chanx_right_in[12], chanx_left_in[18], chanx_right_in[18], chanx_left_in[24], chanx_right_in[24], chanx_left_in[30], chanx_right_in[30], chanx_left_in[36], chanx_right_in[36], chanx_left_in[42], chanx_right_in[42], chanx_left_in[48], chanx_right_in[48], chanx_left_in[54], chanx_right_in[54], chanx_left_in[60], chanx_right_in[60], chanx_left_in[66], chanx_right_in[66], chanx_left_in[72], chanx_right_in[72], chanx_left_in[75], chanx_right_in[75], chanx_left_in[81], chanx_right_in[81], chanx_left_in[87], chanx_right_in[87], chanx_left_in[93], chanx_right_in[93], chanx_left_in[99], chanx_right_in[99], chanx_left_in[105], chanx_right_in[105], chanx_left_in[111], chanx_right_in[111], chanx_left_in[117], chanx_right_in[117], chanx_left_in[123], chanx_right_in[123], chanx_left_in[129], chanx_right_in[129], chanx_left_in[135], chanx_right_in[135], chanx_left_in[141], chanx_right_in[141], chanx_left_in[147], chanx_right_in[147], chanx_left_in[153], chanx_right_in[153], chanx_left_in[159], chanx_right_in[159], chanx_left_in[165], chanx_right_in[165], chanx_left_in[171], chanx_right_in[171], chanx_left_in[177], chanx_right_in[177], chanx_left_in[183], chanx_right_in[183], chanx_left_in[189], chanx_right_in[189], chanx_left_in[195], chanx_right_in[195], chanx_left_in[201], chanx_right_in[201], chanx_left_in[207], chanx_right_in[207], chanx_left_in[213], chanx_right_in[213], chanx_left_in[219], chanx_right_in[219], chanx_left_in[225], chanx_right_in[225], chanx_left_in[231], chanx_right_in[231], chanx_left_in[237], chanx_right_in[237], chanx_left_in[243], chanx_right_in[243], chanx_left_in[249], chanx_right_in[249], chanx_left_in[255], chanx_right_in[255], chanx_left_in[261], chanx_right_in[261], chanx_left_in[267], chanx_right_in[267], chanx_left_in[273], chanx_right_in[273], chanx_left_in[279], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size96_75_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_75_sram_inv[0:6]),
		.out(bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_));

	mux_tree_tapbuf_size96 mux_top_ipin_2 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[7], chanx_right_in[7], chanx_left_in[13], chanx_right_in[13], chanx_left_in[19], chanx_right_in[19], chanx_left_in[25], chanx_right_in[25], chanx_left_in[31], chanx_right_in[31], chanx_left_in[37], chanx_right_in[37], chanx_left_in[43], chanx_right_in[43], chanx_left_in[49], chanx_right_in[49], chanx_left_in[55], chanx_right_in[55], chanx_left_in[61], chanx_right_in[61], chanx_left_in[67], chanx_right_in[67], chanx_left_in[73], chanx_right_in[73], chanx_left_in[76], chanx_right_in[76], chanx_left_in[82], chanx_right_in[82], chanx_left_in[88], chanx_right_in[88], chanx_left_in[94], chanx_right_in[94], chanx_left_in[100], chanx_right_in[100], chanx_left_in[106], chanx_right_in[106], chanx_left_in[112], chanx_right_in[112], chanx_left_in[118], chanx_right_in[118], chanx_left_in[124], chanx_right_in[124], chanx_left_in[130], chanx_right_in[130], chanx_left_in[136], chanx_right_in[136], chanx_left_in[142], chanx_right_in[142], chanx_left_in[148], chanx_right_in[148], chanx_left_in[154], chanx_right_in[154], chanx_left_in[160], chanx_right_in[160], chanx_left_in[166], chanx_right_in[166], chanx_left_in[172], chanx_right_in[172], chanx_left_in[178], chanx_right_in[178], chanx_left_in[184], chanx_right_in[184], chanx_left_in[190], chanx_right_in[190], chanx_left_in[196], chanx_right_in[196], chanx_left_in[202], chanx_right_in[202], chanx_left_in[208], chanx_right_in[208], chanx_left_in[214], chanx_right_in[214], chanx_left_in[220], chanx_right_in[220], chanx_left_in[226], chanx_right_in[226], chanx_left_in[232], chanx_right_in[232], chanx_left_in[238], chanx_right_in[238], chanx_left_in[244], chanx_right_in[244], chanx_left_in[250], chanx_right_in[250], chanx_left_in[256], chanx_right_in[256], chanx_left_in[262], chanx_right_in[262], chanx_left_in[268], chanx_right_in[268], chanx_left_in[274], chanx_right_in[274], chanx_left_in[280], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size96_76_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size96_76_sram_inv[0:6]),
		.out(bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size96_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_0_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_0_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_1_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_1_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_2_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_2_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_3_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_3_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_4_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_4_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_5_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_5_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_6_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_6_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_7_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_7_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_8_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_8_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_9_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_9_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_10_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_10_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_11_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_11_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_12_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_12_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_13_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_13_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_14_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_14_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_15_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_15_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_16_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_16_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_17_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_17_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_18_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_18_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_19_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_19_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_20_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_20_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_21_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_21_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_22_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_22_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_23_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_23_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_24_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_24_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_25_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_25_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_26_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_26_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_27_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_27_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_28_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_28_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_29_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_29_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_30_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_30_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_31_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_31_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_32_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_32_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_33_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_33_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_34_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_34_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_35_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_35_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_36_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_36_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_37_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_37_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_38_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_38_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_39_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_39_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_40_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_40_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_41_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_41_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_42_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_42_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_43_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_43_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_44_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_44_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_45_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_45_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_46_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_46_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_47_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_47_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_48_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_48_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_49_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_49_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_50_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_50_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_51_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_51_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_52_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_52_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_53_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_53_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_54_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_54_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_55_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_55_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_56_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_56_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_57_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_57_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_58_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_58_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_59_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_59_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_60_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_60_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_61_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_61_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_62_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_62_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_63_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_63_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_64_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_64_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_65_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_65_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_66_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_66_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_67_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_67_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_68_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_68_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_69_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_69_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_70_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_70_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_71_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_71_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_72_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_72_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_bottom_ipin_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_73_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_73_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_top_ipin_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_74_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_74_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_top_ipin_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size96_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_75_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_75_sram_inv[0:6]));

	mux_tree_tapbuf_size96_mem mem_top_ipin_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size96_mem_75_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size96_76_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size96_76_sram_inv[0:6]));

endmodule
// ----- END Verilog module for cbx_6__5_ -----

//----- Default net type -----
`default_nettype wire




