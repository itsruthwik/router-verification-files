//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][6]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Jun 27 10:27:38 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__6_ -----
module sb_0__6_(prog_clk,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:188] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:188] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:188] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:188] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_100_sram;
wire [0:1] mux_tree_tapbuf_size2_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_101_sram;
wire [0:1] mux_tree_tapbuf_size2_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_102_sram;
wire [0:1] mux_tree_tapbuf_size2_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_103_sram;
wire [0:1] mux_tree_tapbuf_size2_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_104_sram;
wire [0:1] mux_tree_tapbuf_size2_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_105_sram;
wire [0:1] mux_tree_tapbuf_size2_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_106_sram;
wire [0:1] mux_tree_tapbuf_size2_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_107_sram;
wire [0:1] mux_tree_tapbuf_size2_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_108_sram;
wire [0:1] mux_tree_tapbuf_size2_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_109_sram;
wire [0:1] mux_tree_tapbuf_size2_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_110_sram;
wire [0:1] mux_tree_tapbuf_size2_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_111_sram;
wire [0:1] mux_tree_tapbuf_size2_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_112_sram;
wire [0:1] mux_tree_tapbuf_size2_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_113_sram;
wire [0:1] mux_tree_tapbuf_size2_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_114_sram;
wire [0:1] mux_tree_tapbuf_size2_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_115_sram;
wire [0:1] mux_tree_tapbuf_size2_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_116_sram;
wire [0:1] mux_tree_tapbuf_size2_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_117_sram;
wire [0:1] mux_tree_tapbuf_size2_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_118_sram;
wire [0:1] mux_tree_tapbuf_size2_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_119_sram;
wire [0:1] mux_tree_tapbuf_size2_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_120_sram;
wire [0:1] mux_tree_tapbuf_size2_120_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_121_sram;
wire [0:1] mux_tree_tapbuf_size2_121_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_122_sram;
wire [0:1] mux_tree_tapbuf_size2_122_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_123_sram;
wire [0:1] mux_tree_tapbuf_size2_123_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_124_sram;
wire [0:1] mux_tree_tapbuf_size2_124_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_125_sram;
wire [0:1] mux_tree_tapbuf_size2_125_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_126_sram;
wire [0:1] mux_tree_tapbuf_size2_126_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_127_sram;
wire [0:1] mux_tree_tapbuf_size2_127_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_128_sram;
wire [0:1] mux_tree_tapbuf_size2_128_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_129_sram;
wire [0:1] mux_tree_tapbuf_size2_129_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_130_sram;
wire [0:1] mux_tree_tapbuf_size2_130_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_131_sram;
wire [0:1] mux_tree_tapbuf_size2_131_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_132_sram;
wire [0:1] mux_tree_tapbuf_size2_132_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_133_sram;
wire [0:1] mux_tree_tapbuf_size2_133_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_134_sram;
wire [0:1] mux_tree_tapbuf_size2_134_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_135_sram;
wire [0:1] mux_tree_tapbuf_size2_135_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_136_sram;
wire [0:1] mux_tree_tapbuf_size2_136_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_137_sram;
wire [0:1] mux_tree_tapbuf_size2_137_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_138_sram;
wire [0:1] mux_tree_tapbuf_size2_138_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_139_sram;
wire [0:1] mux_tree_tapbuf_size2_139_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_140_sram;
wire [0:1] mux_tree_tapbuf_size2_140_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_141_sram;
wire [0:1] mux_tree_tapbuf_size2_141_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_142_sram;
wire [0:1] mux_tree_tapbuf_size2_142_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_143_sram;
wire [0:1] mux_tree_tapbuf_size2_143_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_144_sram;
wire [0:1] mux_tree_tapbuf_size2_144_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_145_sram;
wire [0:1] mux_tree_tapbuf_size2_145_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_146_sram;
wire [0:1] mux_tree_tapbuf_size2_146_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_147_sram;
wire [0:1] mux_tree_tapbuf_size2_147_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_148_sram;
wire [0:1] mux_tree_tapbuf_size2_148_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_149_sram;
wire [0:1] mux_tree_tapbuf_size2_149_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_150_sram;
wire [0:1] mux_tree_tapbuf_size2_150_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_151_sram;
wire [0:1] mux_tree_tapbuf_size2_151_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_152_sram;
wire [0:1] mux_tree_tapbuf_size2_152_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_153_sram;
wire [0:1] mux_tree_tapbuf_size2_153_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_154_sram;
wire [0:1] mux_tree_tapbuf_size2_154_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_155_sram;
wire [0:1] mux_tree_tapbuf_size2_155_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_156_sram;
wire [0:1] mux_tree_tapbuf_size2_156_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_157_sram;
wire [0:1] mux_tree_tapbuf_size2_157_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_158_sram;
wire [0:1] mux_tree_tapbuf_size2_158_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_159_sram;
wire [0:1] mux_tree_tapbuf_size2_159_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_160_sram;
wire [0:1] mux_tree_tapbuf_size2_160_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_161_sram;
wire [0:1] mux_tree_tapbuf_size2_161_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_162_sram;
wire [0:1] mux_tree_tapbuf_size2_162_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_163_sram;
wire [0:1] mux_tree_tapbuf_size2_163_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_164_sram;
wire [0:1] mux_tree_tapbuf_size2_164_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_165_sram;
wire [0:1] mux_tree_tapbuf_size2_165_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_166_sram;
wire [0:1] mux_tree_tapbuf_size2_166_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_167_sram;
wire [0:1] mux_tree_tapbuf_size2_167_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_168_sram;
wire [0:1] mux_tree_tapbuf_size2_168_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_169_sram;
wire [0:1] mux_tree_tapbuf_size2_169_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_16_sram;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_170_sram;
wire [0:1] mux_tree_tapbuf_size2_170_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_171_sram;
wire [0:1] mux_tree_tapbuf_size2_171_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_172_sram;
wire [0:1] mux_tree_tapbuf_size2_172_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_173_sram;
wire [0:1] mux_tree_tapbuf_size2_173_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_174_sram;
wire [0:1] mux_tree_tapbuf_size2_174_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_175_sram;
wire [0:1] mux_tree_tapbuf_size2_175_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_176_sram;
wire [0:1] mux_tree_tapbuf_size2_176_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_177_sram;
wire [0:1] mux_tree_tapbuf_size2_177_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_178_sram;
wire [0:1] mux_tree_tapbuf_size2_178_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_179_sram;
wire [0:1] mux_tree_tapbuf_size2_179_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_17_sram;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_180_sram;
wire [0:1] mux_tree_tapbuf_size2_180_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_181_sram;
wire [0:1] mux_tree_tapbuf_size2_181_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_182_sram;
wire [0:1] mux_tree_tapbuf_size2_182_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_183_sram;
wire [0:1] mux_tree_tapbuf_size2_183_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_184_sram;
wire [0:1] mux_tree_tapbuf_size2_184_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_185_sram;
wire [0:1] mux_tree_tapbuf_size2_185_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_186_sram;
wire [0:1] mux_tree_tapbuf_size2_186_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_187_sram;
wire [0:1] mux_tree_tapbuf_size2_187_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_188_sram;
wire [0:1] mux_tree_tapbuf_size2_188_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_189_sram;
wire [0:1] mux_tree_tapbuf_size2_189_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_18_sram;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_190_sram;
wire [0:1] mux_tree_tapbuf_size2_190_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_191_sram;
wire [0:1] mux_tree_tapbuf_size2_191_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_192_sram;
wire [0:1] mux_tree_tapbuf_size2_192_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_193_sram;
wire [0:1] mux_tree_tapbuf_size2_193_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_194_sram;
wire [0:1] mux_tree_tapbuf_size2_194_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_195_sram;
wire [0:1] mux_tree_tapbuf_size2_195_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_196_sram;
wire [0:1] mux_tree_tapbuf_size2_196_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_197_sram;
wire [0:1] mux_tree_tapbuf_size2_197_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_198_sram;
wire [0:1] mux_tree_tapbuf_size2_198_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_199_sram;
wire [0:1] mux_tree_tapbuf_size2_199_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_19_sram;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_200_sram;
wire [0:1] mux_tree_tapbuf_size2_200_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_201_sram;
wire [0:1] mux_tree_tapbuf_size2_201_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_202_sram;
wire [0:1] mux_tree_tapbuf_size2_202_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_203_sram;
wire [0:1] mux_tree_tapbuf_size2_203_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_204_sram;
wire [0:1] mux_tree_tapbuf_size2_204_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_205_sram;
wire [0:1] mux_tree_tapbuf_size2_205_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_206_sram;
wire [0:1] mux_tree_tapbuf_size2_206_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_207_sram;
wire [0:1] mux_tree_tapbuf_size2_207_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_208_sram;
wire [0:1] mux_tree_tapbuf_size2_208_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_209_sram;
wire [0:1] mux_tree_tapbuf_size2_209_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_20_sram;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_210_sram;
wire [0:1] mux_tree_tapbuf_size2_210_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_211_sram;
wire [0:1] mux_tree_tapbuf_size2_211_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_212_sram;
wire [0:1] mux_tree_tapbuf_size2_212_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_213_sram;
wire [0:1] mux_tree_tapbuf_size2_213_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_214_sram;
wire [0:1] mux_tree_tapbuf_size2_214_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_215_sram;
wire [0:1] mux_tree_tapbuf_size2_215_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_216_sram;
wire [0:1] mux_tree_tapbuf_size2_216_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_217_sram;
wire [0:1] mux_tree_tapbuf_size2_217_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_218_sram;
wire [0:1] mux_tree_tapbuf_size2_218_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_219_sram;
wire [0:1] mux_tree_tapbuf_size2_219_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_21_sram;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_220_sram;
wire [0:1] mux_tree_tapbuf_size2_220_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_221_sram;
wire [0:1] mux_tree_tapbuf_size2_221_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_222_sram;
wire [0:1] mux_tree_tapbuf_size2_222_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_223_sram;
wire [0:1] mux_tree_tapbuf_size2_223_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_224_sram;
wire [0:1] mux_tree_tapbuf_size2_224_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_225_sram;
wire [0:1] mux_tree_tapbuf_size2_225_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_226_sram;
wire [0:1] mux_tree_tapbuf_size2_226_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_227_sram;
wire [0:1] mux_tree_tapbuf_size2_227_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_228_sram;
wire [0:1] mux_tree_tapbuf_size2_228_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_229_sram;
wire [0:1] mux_tree_tapbuf_size2_229_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_22_sram;
wire [0:1] mux_tree_tapbuf_size2_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_230_sram;
wire [0:1] mux_tree_tapbuf_size2_230_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_231_sram;
wire [0:1] mux_tree_tapbuf_size2_231_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_232_sram;
wire [0:1] mux_tree_tapbuf_size2_232_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_233_sram;
wire [0:1] mux_tree_tapbuf_size2_233_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_234_sram;
wire [0:1] mux_tree_tapbuf_size2_234_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_235_sram;
wire [0:1] mux_tree_tapbuf_size2_235_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_236_sram;
wire [0:1] mux_tree_tapbuf_size2_236_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_237_sram;
wire [0:1] mux_tree_tapbuf_size2_237_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_238_sram;
wire [0:1] mux_tree_tapbuf_size2_238_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_239_sram;
wire [0:1] mux_tree_tapbuf_size2_239_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_23_sram;
wire [0:1] mux_tree_tapbuf_size2_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_240_sram;
wire [0:1] mux_tree_tapbuf_size2_240_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_241_sram;
wire [0:1] mux_tree_tapbuf_size2_241_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_242_sram;
wire [0:1] mux_tree_tapbuf_size2_242_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_243_sram;
wire [0:1] mux_tree_tapbuf_size2_243_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_244_sram;
wire [0:1] mux_tree_tapbuf_size2_244_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_245_sram;
wire [0:1] mux_tree_tapbuf_size2_245_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_246_sram;
wire [0:1] mux_tree_tapbuf_size2_246_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_247_sram;
wire [0:1] mux_tree_tapbuf_size2_247_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_248_sram;
wire [0:1] mux_tree_tapbuf_size2_248_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_249_sram;
wire [0:1] mux_tree_tapbuf_size2_249_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_24_sram;
wire [0:1] mux_tree_tapbuf_size2_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_250_sram;
wire [0:1] mux_tree_tapbuf_size2_250_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_251_sram;
wire [0:1] mux_tree_tapbuf_size2_251_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_252_sram;
wire [0:1] mux_tree_tapbuf_size2_252_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_253_sram;
wire [0:1] mux_tree_tapbuf_size2_253_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_254_sram;
wire [0:1] mux_tree_tapbuf_size2_254_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_255_sram;
wire [0:1] mux_tree_tapbuf_size2_255_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_256_sram;
wire [0:1] mux_tree_tapbuf_size2_256_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_257_sram;
wire [0:1] mux_tree_tapbuf_size2_257_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_258_sram;
wire [0:1] mux_tree_tapbuf_size2_258_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_259_sram;
wire [0:1] mux_tree_tapbuf_size2_259_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_25_sram;
wire [0:1] mux_tree_tapbuf_size2_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_260_sram;
wire [0:1] mux_tree_tapbuf_size2_260_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_261_sram;
wire [0:1] mux_tree_tapbuf_size2_261_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_262_sram;
wire [0:1] mux_tree_tapbuf_size2_262_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_263_sram;
wire [0:1] mux_tree_tapbuf_size2_263_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_264_sram;
wire [0:1] mux_tree_tapbuf_size2_264_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_265_sram;
wire [0:1] mux_tree_tapbuf_size2_265_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_266_sram;
wire [0:1] mux_tree_tapbuf_size2_266_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_267_sram;
wire [0:1] mux_tree_tapbuf_size2_267_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_268_sram;
wire [0:1] mux_tree_tapbuf_size2_268_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_269_sram;
wire [0:1] mux_tree_tapbuf_size2_269_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_26_sram;
wire [0:1] mux_tree_tapbuf_size2_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_270_sram;
wire [0:1] mux_tree_tapbuf_size2_270_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_271_sram;
wire [0:1] mux_tree_tapbuf_size2_271_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_272_sram;
wire [0:1] mux_tree_tapbuf_size2_272_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_273_sram;
wire [0:1] mux_tree_tapbuf_size2_273_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_274_sram;
wire [0:1] mux_tree_tapbuf_size2_274_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_275_sram;
wire [0:1] mux_tree_tapbuf_size2_275_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_276_sram;
wire [0:1] mux_tree_tapbuf_size2_276_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_277_sram;
wire [0:1] mux_tree_tapbuf_size2_277_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_278_sram;
wire [0:1] mux_tree_tapbuf_size2_278_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_279_sram;
wire [0:1] mux_tree_tapbuf_size2_279_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_27_sram;
wire [0:1] mux_tree_tapbuf_size2_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_280_sram;
wire [0:1] mux_tree_tapbuf_size2_280_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_281_sram;
wire [0:1] mux_tree_tapbuf_size2_281_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_282_sram;
wire [0:1] mux_tree_tapbuf_size2_282_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_283_sram;
wire [0:1] mux_tree_tapbuf_size2_283_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_284_sram;
wire [0:1] mux_tree_tapbuf_size2_284_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_285_sram;
wire [0:1] mux_tree_tapbuf_size2_285_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_286_sram;
wire [0:1] mux_tree_tapbuf_size2_286_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_287_sram;
wire [0:1] mux_tree_tapbuf_size2_287_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_288_sram;
wire [0:1] mux_tree_tapbuf_size2_288_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_289_sram;
wire [0:1] mux_tree_tapbuf_size2_289_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_28_sram;
wire [0:1] mux_tree_tapbuf_size2_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_290_sram;
wire [0:1] mux_tree_tapbuf_size2_290_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_291_sram;
wire [0:1] mux_tree_tapbuf_size2_291_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_292_sram;
wire [0:1] mux_tree_tapbuf_size2_292_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_293_sram;
wire [0:1] mux_tree_tapbuf_size2_293_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_294_sram;
wire [0:1] mux_tree_tapbuf_size2_294_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_295_sram;
wire [0:1] mux_tree_tapbuf_size2_295_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_296_sram;
wire [0:1] mux_tree_tapbuf_size2_296_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_297_sram;
wire [0:1] mux_tree_tapbuf_size2_297_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_298_sram;
wire [0:1] mux_tree_tapbuf_size2_298_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_299_sram;
wire [0:1] mux_tree_tapbuf_size2_299_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_29_sram;
wire [0:1] mux_tree_tapbuf_size2_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_300_sram;
wire [0:1] mux_tree_tapbuf_size2_300_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_301_sram;
wire [0:1] mux_tree_tapbuf_size2_301_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_302_sram;
wire [0:1] mux_tree_tapbuf_size2_302_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_303_sram;
wire [0:1] mux_tree_tapbuf_size2_303_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_304_sram;
wire [0:1] mux_tree_tapbuf_size2_304_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_305_sram;
wire [0:1] mux_tree_tapbuf_size2_305_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_306_sram;
wire [0:1] mux_tree_tapbuf_size2_306_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_307_sram;
wire [0:1] mux_tree_tapbuf_size2_307_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_308_sram;
wire [0:1] mux_tree_tapbuf_size2_308_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_309_sram;
wire [0:1] mux_tree_tapbuf_size2_309_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_30_sram;
wire [0:1] mux_tree_tapbuf_size2_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_310_sram;
wire [0:1] mux_tree_tapbuf_size2_310_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_311_sram;
wire [0:1] mux_tree_tapbuf_size2_311_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_312_sram;
wire [0:1] mux_tree_tapbuf_size2_312_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_313_sram;
wire [0:1] mux_tree_tapbuf_size2_313_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_314_sram;
wire [0:1] mux_tree_tapbuf_size2_314_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_315_sram;
wire [0:1] mux_tree_tapbuf_size2_315_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_316_sram;
wire [0:1] mux_tree_tapbuf_size2_316_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_317_sram;
wire [0:1] mux_tree_tapbuf_size2_317_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_318_sram;
wire [0:1] mux_tree_tapbuf_size2_318_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_319_sram;
wire [0:1] mux_tree_tapbuf_size2_319_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_31_sram;
wire [0:1] mux_tree_tapbuf_size2_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_320_sram;
wire [0:1] mux_tree_tapbuf_size2_320_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_321_sram;
wire [0:1] mux_tree_tapbuf_size2_321_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_322_sram;
wire [0:1] mux_tree_tapbuf_size2_322_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_323_sram;
wire [0:1] mux_tree_tapbuf_size2_323_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_324_sram;
wire [0:1] mux_tree_tapbuf_size2_324_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_325_sram;
wire [0:1] mux_tree_tapbuf_size2_325_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_326_sram;
wire [0:1] mux_tree_tapbuf_size2_326_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_327_sram;
wire [0:1] mux_tree_tapbuf_size2_327_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_328_sram;
wire [0:1] mux_tree_tapbuf_size2_328_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_329_sram;
wire [0:1] mux_tree_tapbuf_size2_329_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_32_sram;
wire [0:1] mux_tree_tapbuf_size2_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_330_sram;
wire [0:1] mux_tree_tapbuf_size2_330_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_331_sram;
wire [0:1] mux_tree_tapbuf_size2_331_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_332_sram;
wire [0:1] mux_tree_tapbuf_size2_332_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_333_sram;
wire [0:1] mux_tree_tapbuf_size2_333_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_334_sram;
wire [0:1] mux_tree_tapbuf_size2_334_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_335_sram;
wire [0:1] mux_tree_tapbuf_size2_335_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_336_sram;
wire [0:1] mux_tree_tapbuf_size2_336_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_337_sram;
wire [0:1] mux_tree_tapbuf_size2_337_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_338_sram;
wire [0:1] mux_tree_tapbuf_size2_338_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_339_sram;
wire [0:1] mux_tree_tapbuf_size2_339_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_33_sram;
wire [0:1] mux_tree_tapbuf_size2_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_340_sram;
wire [0:1] mux_tree_tapbuf_size2_340_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_341_sram;
wire [0:1] mux_tree_tapbuf_size2_341_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_342_sram;
wire [0:1] mux_tree_tapbuf_size2_342_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_343_sram;
wire [0:1] mux_tree_tapbuf_size2_343_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_344_sram;
wire [0:1] mux_tree_tapbuf_size2_344_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_345_sram;
wire [0:1] mux_tree_tapbuf_size2_345_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_346_sram;
wire [0:1] mux_tree_tapbuf_size2_346_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_347_sram;
wire [0:1] mux_tree_tapbuf_size2_347_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_348_sram;
wire [0:1] mux_tree_tapbuf_size2_348_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_349_sram;
wire [0:1] mux_tree_tapbuf_size2_349_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_34_sram;
wire [0:1] mux_tree_tapbuf_size2_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_350_sram;
wire [0:1] mux_tree_tapbuf_size2_350_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_351_sram;
wire [0:1] mux_tree_tapbuf_size2_351_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_352_sram;
wire [0:1] mux_tree_tapbuf_size2_352_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_353_sram;
wire [0:1] mux_tree_tapbuf_size2_353_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_354_sram;
wire [0:1] mux_tree_tapbuf_size2_354_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_355_sram;
wire [0:1] mux_tree_tapbuf_size2_355_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_356_sram;
wire [0:1] mux_tree_tapbuf_size2_356_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_357_sram;
wire [0:1] mux_tree_tapbuf_size2_357_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_358_sram;
wire [0:1] mux_tree_tapbuf_size2_358_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_359_sram;
wire [0:1] mux_tree_tapbuf_size2_359_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_35_sram;
wire [0:1] mux_tree_tapbuf_size2_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_360_sram;
wire [0:1] mux_tree_tapbuf_size2_360_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_361_sram;
wire [0:1] mux_tree_tapbuf_size2_361_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_362_sram;
wire [0:1] mux_tree_tapbuf_size2_362_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_363_sram;
wire [0:1] mux_tree_tapbuf_size2_363_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_364_sram;
wire [0:1] mux_tree_tapbuf_size2_364_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_365_sram;
wire [0:1] mux_tree_tapbuf_size2_365_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_366_sram;
wire [0:1] mux_tree_tapbuf_size2_366_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_367_sram;
wire [0:1] mux_tree_tapbuf_size2_367_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_368_sram;
wire [0:1] mux_tree_tapbuf_size2_368_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_369_sram;
wire [0:1] mux_tree_tapbuf_size2_369_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_36_sram;
wire [0:1] mux_tree_tapbuf_size2_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_370_sram;
wire [0:1] mux_tree_tapbuf_size2_370_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_371_sram;
wire [0:1] mux_tree_tapbuf_size2_371_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_372_sram;
wire [0:1] mux_tree_tapbuf_size2_372_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_373_sram;
wire [0:1] mux_tree_tapbuf_size2_373_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_374_sram;
wire [0:1] mux_tree_tapbuf_size2_374_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_375_sram;
wire [0:1] mux_tree_tapbuf_size2_375_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_376_sram;
wire [0:1] mux_tree_tapbuf_size2_376_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_377_sram;
wire [0:1] mux_tree_tapbuf_size2_377_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_37_sram;
wire [0:1] mux_tree_tapbuf_size2_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_38_sram;
wire [0:1] mux_tree_tapbuf_size2_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_39_sram;
wire [0:1] mux_tree_tapbuf_size2_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_40_sram;
wire [0:1] mux_tree_tapbuf_size2_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_41_sram;
wire [0:1] mux_tree_tapbuf_size2_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_42_sram;
wire [0:1] mux_tree_tapbuf_size2_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_43_sram;
wire [0:1] mux_tree_tapbuf_size2_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_44_sram;
wire [0:1] mux_tree_tapbuf_size2_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_45_sram;
wire [0:1] mux_tree_tapbuf_size2_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_46_sram;
wire [0:1] mux_tree_tapbuf_size2_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_47_sram;
wire [0:1] mux_tree_tapbuf_size2_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_48_sram;
wire [0:1] mux_tree_tapbuf_size2_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_49_sram;
wire [0:1] mux_tree_tapbuf_size2_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_50_sram;
wire [0:1] mux_tree_tapbuf_size2_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_51_sram;
wire [0:1] mux_tree_tapbuf_size2_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_52_sram;
wire [0:1] mux_tree_tapbuf_size2_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_53_sram;
wire [0:1] mux_tree_tapbuf_size2_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_54_sram;
wire [0:1] mux_tree_tapbuf_size2_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_55_sram;
wire [0:1] mux_tree_tapbuf_size2_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_56_sram;
wire [0:1] mux_tree_tapbuf_size2_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_57_sram;
wire [0:1] mux_tree_tapbuf_size2_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_58_sram;
wire [0:1] mux_tree_tapbuf_size2_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_59_sram;
wire [0:1] mux_tree_tapbuf_size2_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_60_sram;
wire [0:1] mux_tree_tapbuf_size2_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_61_sram;
wire [0:1] mux_tree_tapbuf_size2_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_62_sram;
wire [0:1] mux_tree_tapbuf_size2_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_63_sram;
wire [0:1] mux_tree_tapbuf_size2_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_64_sram;
wire [0:1] mux_tree_tapbuf_size2_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_65_sram;
wire [0:1] mux_tree_tapbuf_size2_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_66_sram;
wire [0:1] mux_tree_tapbuf_size2_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_67_sram;
wire [0:1] mux_tree_tapbuf_size2_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_68_sram;
wire [0:1] mux_tree_tapbuf_size2_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_69_sram;
wire [0:1] mux_tree_tapbuf_size2_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_70_sram;
wire [0:1] mux_tree_tapbuf_size2_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_71_sram;
wire [0:1] mux_tree_tapbuf_size2_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_72_sram;
wire [0:1] mux_tree_tapbuf_size2_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_73_sram;
wire [0:1] mux_tree_tapbuf_size2_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_74_sram;
wire [0:1] mux_tree_tapbuf_size2_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_75_sram;
wire [0:1] mux_tree_tapbuf_size2_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_76_sram;
wire [0:1] mux_tree_tapbuf_size2_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_77_sram;
wire [0:1] mux_tree_tapbuf_size2_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_78_sram;
wire [0:1] mux_tree_tapbuf_size2_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_79_sram;
wire [0:1] mux_tree_tapbuf_size2_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_80_sram;
wire [0:1] mux_tree_tapbuf_size2_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_81_sram;
wire [0:1] mux_tree_tapbuf_size2_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_82_sram;
wire [0:1] mux_tree_tapbuf_size2_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_83_sram;
wire [0:1] mux_tree_tapbuf_size2_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_84_sram;
wire [0:1] mux_tree_tapbuf_size2_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_85_sram;
wire [0:1] mux_tree_tapbuf_size2_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_86_sram;
wire [0:1] mux_tree_tapbuf_size2_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_87_sram;
wire [0:1] mux_tree_tapbuf_size2_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_88_sram;
wire [0:1] mux_tree_tapbuf_size2_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_89_sram;
wire [0:1] mux_tree_tapbuf_size2_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_90_sram;
wire [0:1] mux_tree_tapbuf_size2_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_91_sram;
wire [0:1] mux_tree_tapbuf_size2_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_92_sram;
wire [0:1] mux_tree_tapbuf_size2_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_93_sram;
wire [0:1] mux_tree_tapbuf_size2_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_94_sram;
wire [0:1] mux_tree_tapbuf_size2_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_95_sram;
wire [0:1] mux_tree_tapbuf_size2_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_96_sram;
wire [0:1] mux_tree_tapbuf_size2_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_97_sram;
wire [0:1] mux_tree_tapbuf_size2_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_98_sram;
wire [0:1] mux_tree_tapbuf_size2_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_99_sram;
wire [0:1] mux_tree_tapbuf_size2_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_136_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_137_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_138_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_139_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_140_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_141_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_142_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_143_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_144_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_145_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_146_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_147_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_148_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_149_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_150_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_151_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_152_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_153_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_154_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_155_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_156_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_157_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_158_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_159_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_160_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_161_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_162_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_163_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_164_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_165_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_166_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_167_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_168_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_169_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_170_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_171_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_172_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_173_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_174_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_175_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_176_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_177_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_178_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_179_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_180_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_181_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_182_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_183_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_184_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_185_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_186_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_187_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_188_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_189_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_190_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_191_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_192_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_193_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_194_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_195_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_196_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_197_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_198_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_199_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_200_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_201_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_202_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_203_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_204_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_205_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_206_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_207_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_208_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_209_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_210_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_211_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_212_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_213_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_214_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_215_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_216_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_217_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_218_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_219_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_220_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_221_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_222_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_223_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_224_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_225_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_226_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_227_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_228_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_229_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_230_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_231_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_232_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_233_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_234_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_235_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_236_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_237_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_238_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_239_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_240_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_241_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_242_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_243_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_244_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_245_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_246_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_247_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_248_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_249_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_250_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_251_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_252_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_253_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_254_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_255_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_256_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_257_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_258_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_259_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_260_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_261_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_262_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_263_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_264_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_265_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_266_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_267_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_268_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_269_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_270_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_271_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_272_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_273_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_274_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_275_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_276_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_277_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_278_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_279_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_280_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_281_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_282_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_283_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_284_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_285_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_286_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_287_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_288_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_289_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_290_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_291_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_292_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_293_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_294_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_295_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_296_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_297_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_298_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_299_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_300_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_301_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_302_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_303_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_304_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_305_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_306_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_307_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_308_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_309_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_310_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_311_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_312_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_313_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_314_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_315_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_316_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_317_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_318_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_319_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_320_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_321_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_322_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_323_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_324_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_325_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_326_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_327_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_328_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_329_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_330_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_331_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_332_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_333_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_334_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_335_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_336_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_337_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_338_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_339_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_340_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_341_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_342_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_343_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_344_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_345_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_346_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_347_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_348_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_349_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_350_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_351_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_352_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_353_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_354_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_355_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_356_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_357_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_358_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_359_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_360_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_361_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_362_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_363_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_364_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_365_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_366_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_367_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_368_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_369_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_370_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_371_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_372_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_373_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_374_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_375_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_376_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size2 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[187]}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size2 mux_right_track_2 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[186]}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_size2 mux_right_track_4 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[185]}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_size2 mux_right_track_6 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[184]}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_size2 mux_right_track_8 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[183]}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size2 mux_right_track_10 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[182]}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_size2 mux_right_track_12 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[181]}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_size2 mux_right_track_14 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[180]}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_size2 mux_right_track_16 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[179]}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size2 mux_right_track_18 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[178]}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_size2 mux_right_track_20 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[177]}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_size2 mux_right_track_22 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[176]}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_size2 mux_right_track_24 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[175]}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size2 mux_right_track_26 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[174]}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_size2 mux_right_track_28 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[173]}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_size2 mux_right_track_30 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[172]}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_size2 mux_right_track_32 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[171]}),
		.sram(mux_tree_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_16_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size2 mux_right_track_34 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[170]}),
		.sram(mux_tree_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_17_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_size2 mux_right_track_36 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[169]}),
		.sram(mux_tree_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_18_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_size2 mux_right_track_38 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[168]}),
		.sram(mux_tree_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_19_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_size2 mux_right_track_40 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[167]}),
		.sram(mux_tree_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_20_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size2 mux_right_track_42 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[166]}),
		.sram(mux_tree_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_21_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_tree_tapbuf_size2 mux_right_track_44 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[165]}),
		.sram(mux_tree_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_22_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_size2 mux_right_track_46 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[164]}),
		.sram(mux_tree_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_23_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_size2 mux_right_track_48 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[163]}),
		.sram(mux_tree_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_24_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size2 mux_right_track_50 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[162]}),
		.sram(mux_tree_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_25_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_tree_tapbuf_size2 mux_right_track_52 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[161]}),
		.sram(mux_tree_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_26_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_size2 mux_right_track_54 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[160]}),
		.sram(mux_tree_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_27_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_size2 mux_right_track_56 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[159]}),
		.sram(mux_tree_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_28_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size2 mux_right_track_58 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[158]}),
		.sram(mux_tree_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_29_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_tree_tapbuf_size2 mux_right_track_60 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[157]}),
		.sram(mux_tree_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_30_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_size2 mux_right_track_62 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[156]}),
		.sram(mux_tree_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_31_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_size2 mux_right_track_64 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[155]}),
		.sram(mux_tree_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_32_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size2 mux_right_track_66 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[154]}),
		.sram(mux_tree_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_33_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_tree_tapbuf_size2 mux_right_track_68 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[153]}),
		.sram(mux_tree_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_34_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_size2 mux_right_track_70 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[152]}),
		.sram(mux_tree_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_35_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_size2 mux_right_track_72 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[151]}),
		.sram(mux_tree_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_36_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size2 mux_right_track_74 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[150]}),
		.sram(mux_tree_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_37_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_tree_tapbuf_size2 mux_right_track_76 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[149]}),
		.sram(mux_tree_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_38_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_size2 mux_right_track_78 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[148]}),
		.sram(mux_tree_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_39_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_size2 mux_right_track_80 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[147]}),
		.sram(mux_tree_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_40_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size2 mux_right_track_82 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[146]}),
		.sram(mux_tree_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_41_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_tree_tapbuf_size2 mux_right_track_84 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[145]}),
		.sram(mux_tree_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_42_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_size2 mux_right_track_86 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[144]}),
		.sram(mux_tree_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_43_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_size2 mux_right_track_88 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[143]}),
		.sram(mux_tree_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_44_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size2 mux_right_track_90 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[142]}),
		.sram(mux_tree_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_45_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_tree_tapbuf_size2 mux_right_track_92 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[141]}),
		.sram(mux_tree_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_46_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_size2 mux_right_track_94 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[140]}),
		.sram(mux_tree_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_47_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_size2 mux_right_track_96 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[139]}),
		.sram(mux_tree_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_48_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size2 mux_right_track_98 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[138]}),
		.sram(mux_tree_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_49_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_tree_tapbuf_size2 mux_right_track_100 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[137]}),
		.sram(mux_tree_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_50_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_size2 mux_right_track_102 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[136]}),
		.sram(mux_tree_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_51_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_size2 mux_right_track_104 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[135]}),
		.sram(mux_tree_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_52_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size2 mux_right_track_106 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[134]}),
		.sram(mux_tree_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_53_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	mux_tree_tapbuf_size2 mux_right_track_108 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[133]}),
		.sram(mux_tree_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_54_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_size2 mux_right_track_110 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[132]}),
		.sram(mux_tree_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_55_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_size2 mux_right_track_112 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[131]}),
		.sram(mux_tree_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_56_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size2 mux_right_track_114 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[130]}),
		.sram(mux_tree_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_57_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_tree_tapbuf_size2 mux_right_track_116 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[129]}),
		.sram(mux_tree_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_58_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_size2 mux_right_track_118 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[128]}),
		.sram(mux_tree_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_59_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_size2 mux_right_track_120 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[127]}),
		.sram(mux_tree_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_60_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size2 mux_right_track_122 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[126]}),
		.sram(mux_tree_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_61_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_tree_tapbuf_size2 mux_right_track_124 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[125]}),
		.sram(mux_tree_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_62_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_size2 mux_right_track_126 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[124]}),
		.sram(mux_tree_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_63_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_size2 mux_right_track_128 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[123]}),
		.sram(mux_tree_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_64_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size2 mux_right_track_130 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[122]}),
		.sram(mux_tree_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_65_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_tree_tapbuf_size2 mux_right_track_132 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[121]}),
		.sram(mux_tree_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_66_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_tree_tapbuf_size2 mux_right_track_134 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[120]}),
		.sram(mux_tree_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_67_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_size2 mux_right_track_136 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[119]}),
		.sram(mux_tree_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_68_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size2 mux_right_track_138 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[118]}),
		.sram(mux_tree_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_69_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_tree_tapbuf_size2 mux_right_track_140 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[117]}),
		.sram(mux_tree_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_70_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_tree_tapbuf_size2 mux_right_track_142 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[116]}),
		.sram(mux_tree_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_71_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_size2 mux_right_track_144 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[115]}),
		.sram(mux_tree_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_72_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size2 mux_right_track_146 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[114]}),
		.sram(mux_tree_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_73_sram_inv[0:1]),
		.out(chanx_right_out[73]));

	mux_tree_tapbuf_size2 mux_right_track_148 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[113]}),
		.sram(mux_tree_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_74_sram_inv[0:1]),
		.out(chanx_right_out[74]));

	mux_tree_tapbuf_size2 mux_right_track_150 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[112]}),
		.sram(mux_tree_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_75_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_size2 mux_right_track_152 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[111]}),
		.sram(mux_tree_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_76_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size2 mux_right_track_154 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[110]}),
		.sram(mux_tree_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_77_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_tree_tapbuf_size2 mux_right_track_156 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[109]}),
		.sram(mux_tree_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_78_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_tree_tapbuf_size2 mux_right_track_158 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[108]}),
		.sram(mux_tree_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_79_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_size2 mux_right_track_160 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[107]}),
		.sram(mux_tree_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_80_sram_inv[0:1]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size2 mux_right_track_162 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[106]}),
		.sram(mux_tree_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_81_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_tree_tapbuf_size2 mux_right_track_164 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[105]}),
		.sram(mux_tree_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_82_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_tree_tapbuf_size2 mux_right_track_166 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[104]}),
		.sram(mux_tree_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_83_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_size2 mux_right_track_168 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[103]}),
		.sram(mux_tree_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_84_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size2 mux_right_track_170 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[102]}),
		.sram(mux_tree_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_85_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_tree_tapbuf_size2 mux_right_track_172 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[101]}),
		.sram(mux_tree_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_86_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_tree_tapbuf_size2 mux_right_track_174 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[100]}),
		.sram(mux_tree_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_87_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_size2 mux_right_track_176 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[99]}),
		.sram(mux_tree_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_88_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size2 mux_right_track_178 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[98]}),
		.sram(mux_tree_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_89_sram_inv[0:1]),
		.out(chanx_right_out[89]));

	mux_tree_tapbuf_size2 mux_right_track_180 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[97]}),
		.sram(mux_tree_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_90_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_tree_tapbuf_size2 mux_right_track_182 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[96]}),
		.sram(mux_tree_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_91_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_size2 mux_right_track_184 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[95]}),
		.sram(mux_tree_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_92_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size2 mux_right_track_186 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[94]}),
		.sram(mux_tree_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_93_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_tree_tapbuf_size2 mux_right_track_188 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[93]}),
		.sram(mux_tree_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_94_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_tree_tapbuf_size2 mux_right_track_190 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[92]}),
		.sram(mux_tree_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_95_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_size2 mux_right_track_192 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[91]}),
		.sram(mux_tree_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_96_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size2 mux_right_track_194 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[90]}),
		.sram(mux_tree_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_97_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_tree_tapbuf_size2 mux_right_track_196 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[89]}),
		.sram(mux_tree_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_98_sram_inv[0:1]),
		.out(chanx_right_out[98]));

	mux_tree_tapbuf_size2 mux_right_track_198 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[88]}),
		.sram(mux_tree_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_99_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_tree_tapbuf_size2 mux_right_track_200 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[87]}),
		.sram(mux_tree_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_100_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size2 mux_right_track_202 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[86]}),
		.sram(mux_tree_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_101_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_tree_tapbuf_size2 mux_right_track_204 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[85]}),
		.sram(mux_tree_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_102_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_tree_tapbuf_size2 mux_right_track_206 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[84]}),
		.sram(mux_tree_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_103_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_tree_tapbuf_size2 mux_right_track_208 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[83]}),
		.sram(mux_tree_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_104_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size2 mux_right_track_210 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[82]}),
		.sram(mux_tree_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_105_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_tree_tapbuf_size2 mux_right_track_212 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[81]}),
		.sram(mux_tree_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_106_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_tree_tapbuf_size2 mux_right_track_214 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[80]}),
		.sram(mux_tree_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_107_sram_inv[0:1]),
		.out(chanx_right_out[107]));

	mux_tree_tapbuf_size2 mux_right_track_216 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[79]}),
		.sram(mux_tree_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_108_sram_inv[0:1]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size2 mux_right_track_218 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[78]}),
		.sram(mux_tree_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_109_sram_inv[0:1]),
		.out(chanx_right_out[109]));

	mux_tree_tapbuf_size2 mux_right_track_220 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[77]}),
		.sram(mux_tree_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_110_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_tree_tapbuf_size2 mux_right_track_222 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[76]}),
		.sram(mux_tree_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_111_sram_inv[0:1]),
		.out(chanx_right_out[111]));

	mux_tree_tapbuf_size2 mux_right_track_224 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[75]}),
		.sram(mux_tree_tapbuf_size2_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_112_sram_inv[0:1]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size2 mux_right_track_226 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[74]}),
		.sram(mux_tree_tapbuf_size2_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_113_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_tree_tapbuf_size2 mux_right_track_228 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[73]}),
		.sram(mux_tree_tapbuf_size2_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_114_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_tree_tapbuf_size2 mux_right_track_230 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[72]}),
		.sram(mux_tree_tapbuf_size2_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_115_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_tree_tapbuf_size2 mux_right_track_232 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[71]}),
		.sram(mux_tree_tapbuf_size2_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_116_sram_inv[0:1]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size2 mux_right_track_234 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[70]}),
		.sram(mux_tree_tapbuf_size2_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_117_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_tree_tapbuf_size2 mux_right_track_236 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[69]}),
		.sram(mux_tree_tapbuf_size2_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_118_sram_inv[0:1]),
		.out(chanx_right_out[118]));

	mux_tree_tapbuf_size2 mux_right_track_238 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[68]}),
		.sram(mux_tree_tapbuf_size2_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_119_sram_inv[0:1]),
		.out(chanx_right_out[119]));

	mux_tree_tapbuf_size2 mux_right_track_240 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[67]}),
		.sram(mux_tree_tapbuf_size2_120_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_120_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size2 mux_right_track_242 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[66]}),
		.sram(mux_tree_tapbuf_size2_121_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_121_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_tree_tapbuf_size2 mux_right_track_244 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[65]}),
		.sram(mux_tree_tapbuf_size2_122_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_122_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_tree_tapbuf_size2 mux_right_track_246 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[64]}),
		.sram(mux_tree_tapbuf_size2_123_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_123_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_tree_tapbuf_size2 mux_right_track_248 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size2_124_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_124_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size2 mux_right_track_250 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[62]}),
		.sram(mux_tree_tapbuf_size2_125_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_125_sram_inv[0:1]),
		.out(chanx_right_out[125]));

	mux_tree_tapbuf_size2 mux_right_track_252 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[61]}),
		.sram(mux_tree_tapbuf_size2_126_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_126_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_tree_tapbuf_size2 mux_right_track_254 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[60]}),
		.sram(mux_tree_tapbuf_size2_127_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_127_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_tree_tapbuf_size2 mux_right_track_256 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_size2_128_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_128_sram_inv[0:1]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size2 mux_right_track_258 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[58]}),
		.sram(mux_tree_tapbuf_size2_129_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_129_sram_inv[0:1]),
		.out(chanx_right_out[129]));

	mux_tree_tapbuf_size2 mux_right_track_260 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[57]}),
		.sram(mux_tree_tapbuf_size2_130_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_130_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_tree_tapbuf_size2 mux_right_track_262 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[56]}),
		.sram(mux_tree_tapbuf_size2_131_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_131_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_tree_tapbuf_size2 mux_right_track_264 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_size2_132_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_132_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size2 mux_right_track_266 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[54]}),
		.sram(mux_tree_tapbuf_size2_133_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_133_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_tree_tapbuf_size2 mux_right_track_268 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[53]}),
		.sram(mux_tree_tapbuf_size2_134_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_134_sram_inv[0:1]),
		.out(chanx_right_out[134]));

	mux_tree_tapbuf_size2 mux_right_track_270 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[52]}),
		.sram(mux_tree_tapbuf_size2_135_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_135_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_tree_tapbuf_size2 mux_right_track_272 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_size2_136_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_136_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size2 mux_right_track_274 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[50]}),
		.sram(mux_tree_tapbuf_size2_137_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_137_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_tree_tapbuf_size2 mux_right_track_276 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[49]}),
		.sram(mux_tree_tapbuf_size2_138_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_138_sram_inv[0:1]),
		.out(chanx_right_out[138]));

	mux_tree_tapbuf_size2 mux_right_track_278 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[48]}),
		.sram(mux_tree_tapbuf_size2_139_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_139_sram_inv[0:1]),
		.out(chanx_right_out[139]));

	mux_tree_tapbuf_size2 mux_right_track_280 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_size2_140_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_140_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size2 mux_right_track_282 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[46]}),
		.sram(mux_tree_tapbuf_size2_141_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_141_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_tree_tapbuf_size2 mux_right_track_284 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[45]}),
		.sram(mux_tree_tapbuf_size2_142_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_142_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_tree_tapbuf_size2 mux_right_track_286 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[44]}),
		.sram(mux_tree_tapbuf_size2_143_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_143_sram_inv[0:1]),
		.out(chanx_right_out[143]));

	mux_tree_tapbuf_size2 mux_right_track_288 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_size2_144_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_144_sram_inv[0:1]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size2 mux_right_track_290 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[42]}),
		.sram(mux_tree_tapbuf_size2_145_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_145_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_tree_tapbuf_size2 mux_right_track_292 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[41]}),
		.sram(mux_tree_tapbuf_size2_146_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_146_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_tree_tapbuf_size2 mux_right_track_294 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[40]}),
		.sram(mux_tree_tapbuf_size2_147_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_147_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_tree_tapbuf_size2 mux_right_track_296 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_size2_148_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_148_sram_inv[0:1]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size2 mux_right_track_298 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[38]}),
		.sram(mux_tree_tapbuf_size2_149_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_149_sram_inv[0:1]),
		.out(chanx_right_out[149]));

	mux_tree_tapbuf_size2 mux_right_track_300 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[37]}),
		.sram(mux_tree_tapbuf_size2_150_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_150_sram_inv[0:1]),
		.out(chanx_right_out[150]));

	mux_tree_tapbuf_size2 mux_right_track_302 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[36]}),
		.sram(mux_tree_tapbuf_size2_151_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_151_sram_inv[0:1]),
		.out(chanx_right_out[151]));

	mux_tree_tapbuf_size2 mux_right_track_304 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_size2_152_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_152_sram_inv[0:1]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size2 mux_right_track_306 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[34]}),
		.sram(mux_tree_tapbuf_size2_153_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_153_sram_inv[0:1]),
		.out(chanx_right_out[153]));

	mux_tree_tapbuf_size2 mux_right_track_308 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[33]}),
		.sram(mux_tree_tapbuf_size2_154_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_154_sram_inv[0:1]),
		.out(chanx_right_out[154]));

	mux_tree_tapbuf_size2 mux_right_track_310 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[32]}),
		.sram(mux_tree_tapbuf_size2_155_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_155_sram_inv[0:1]),
		.out(chanx_right_out[155]));

	mux_tree_tapbuf_size2 mux_right_track_312 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_size2_156_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_156_sram_inv[0:1]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size2 mux_right_track_314 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[30]}),
		.sram(mux_tree_tapbuf_size2_157_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_157_sram_inv[0:1]),
		.out(chanx_right_out[157]));

	mux_tree_tapbuf_size2 mux_right_track_316 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[29]}),
		.sram(mux_tree_tapbuf_size2_158_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_158_sram_inv[0:1]),
		.out(chanx_right_out[158]));

	mux_tree_tapbuf_size2 mux_right_track_318 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[28]}),
		.sram(mux_tree_tapbuf_size2_159_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_159_sram_inv[0:1]),
		.out(chanx_right_out[159]));

	mux_tree_tapbuf_size2 mux_right_track_320 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[27]}),
		.sram(mux_tree_tapbuf_size2_160_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_160_sram_inv[0:1]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size2 mux_right_track_322 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[26]}),
		.sram(mux_tree_tapbuf_size2_161_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_161_sram_inv[0:1]),
		.out(chanx_right_out[161]));

	mux_tree_tapbuf_size2 mux_right_track_324 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[25]}),
		.sram(mux_tree_tapbuf_size2_162_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_162_sram_inv[0:1]),
		.out(chanx_right_out[162]));

	mux_tree_tapbuf_size2 mux_right_track_326 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[24]}),
		.sram(mux_tree_tapbuf_size2_163_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_163_sram_inv[0:1]),
		.out(chanx_right_out[163]));

	mux_tree_tapbuf_size2 mux_right_track_328 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[23]}),
		.sram(mux_tree_tapbuf_size2_164_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_164_sram_inv[0:1]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size2 mux_right_track_330 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[22]}),
		.sram(mux_tree_tapbuf_size2_165_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_165_sram_inv[0:1]),
		.out(chanx_right_out[165]));

	mux_tree_tapbuf_size2 mux_right_track_332 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[21]}),
		.sram(mux_tree_tapbuf_size2_166_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_166_sram_inv[0:1]),
		.out(chanx_right_out[166]));

	mux_tree_tapbuf_size2 mux_right_track_334 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[20]}),
		.sram(mux_tree_tapbuf_size2_167_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_167_sram_inv[0:1]),
		.out(chanx_right_out[167]));

	mux_tree_tapbuf_size2 mux_right_track_336 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[19]}),
		.sram(mux_tree_tapbuf_size2_168_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_168_sram_inv[0:1]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size2 mux_right_track_338 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[18]}),
		.sram(mux_tree_tapbuf_size2_169_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_169_sram_inv[0:1]),
		.out(chanx_right_out[169]));

	mux_tree_tapbuf_size2 mux_right_track_340 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[17]}),
		.sram(mux_tree_tapbuf_size2_170_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_170_sram_inv[0:1]),
		.out(chanx_right_out[170]));

	mux_tree_tapbuf_size2 mux_right_track_342 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[16]}),
		.sram(mux_tree_tapbuf_size2_171_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_171_sram_inv[0:1]),
		.out(chanx_right_out[171]));

	mux_tree_tapbuf_size2 mux_right_track_344 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[15]}),
		.sram(mux_tree_tapbuf_size2_172_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_172_sram_inv[0:1]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size2 mux_right_track_346 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[14]}),
		.sram(mux_tree_tapbuf_size2_173_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_173_sram_inv[0:1]),
		.out(chanx_right_out[173]));

	mux_tree_tapbuf_size2 mux_right_track_348 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[13]}),
		.sram(mux_tree_tapbuf_size2_174_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_174_sram_inv[0:1]),
		.out(chanx_right_out[174]));

	mux_tree_tapbuf_size2 mux_right_track_350 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[12]}),
		.sram(mux_tree_tapbuf_size2_175_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_175_sram_inv[0:1]),
		.out(chanx_right_out[175]));

	mux_tree_tapbuf_size2 mux_right_track_352 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[11]}),
		.sram(mux_tree_tapbuf_size2_176_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_176_sram_inv[0:1]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size2 mux_right_track_354 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[10]}),
		.sram(mux_tree_tapbuf_size2_177_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_177_sram_inv[0:1]),
		.out(chanx_right_out[177]));

	mux_tree_tapbuf_size2 mux_right_track_356 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[9]}),
		.sram(mux_tree_tapbuf_size2_178_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_178_sram_inv[0:1]),
		.out(chanx_right_out[178]));

	mux_tree_tapbuf_size2 mux_right_track_358 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[8]}),
		.sram(mux_tree_tapbuf_size2_179_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_179_sram_inv[0:1]),
		.out(chanx_right_out[179]));

	mux_tree_tapbuf_size2 mux_right_track_360 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[7]}),
		.sram(mux_tree_tapbuf_size2_180_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_180_sram_inv[0:1]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size2 mux_right_track_362 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[6]}),
		.sram(mux_tree_tapbuf_size2_181_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_181_sram_inv[0:1]),
		.out(chanx_right_out[181]));

	mux_tree_tapbuf_size2 mux_right_track_364 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[5]}),
		.sram(mux_tree_tapbuf_size2_182_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_182_sram_inv[0:1]),
		.out(chanx_right_out[182]));

	mux_tree_tapbuf_size2 mux_right_track_366 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[4]}),
		.sram(mux_tree_tapbuf_size2_183_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_183_sram_inv[0:1]),
		.out(chanx_right_out[183]));

	mux_tree_tapbuf_size2 mux_right_track_368 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[3]}),
		.sram(mux_tree_tapbuf_size2_184_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_184_sram_inv[0:1]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size2 mux_right_track_370 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[2]}),
		.sram(mux_tree_tapbuf_size2_185_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_185_sram_inv[0:1]),
		.out(chanx_right_out[185]));

	mux_tree_tapbuf_size2 mux_right_track_372 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[1]}),
		.sram(mux_tree_tapbuf_size2_186_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_186_sram_inv[0:1]),
		.out(chanx_right_out[186]));

	mux_tree_tapbuf_size2 mux_right_track_374 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[0]}),
		.sram(mux_tree_tapbuf_size2_187_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_187_sram_inv[0:1]),
		.out(chanx_right_out[187]));

	mux_tree_tapbuf_size2 mux_right_track_376 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[188]}),
		.sram(mux_tree_tapbuf_size2_188_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_188_sram_inv[0:1]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size2 mux_bottom_track_1 (
		.in({chanx_right_in[187], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_189_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_189_sram_inv[0:1]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size2 mux_bottom_track_3 (
		.in({chanx_right_in[186], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_190_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_190_sram_inv[0:1]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_size2 mux_bottom_track_5 (
		.in({chanx_right_in[185], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_191_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_191_sram_inv[0:1]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_size2 mux_bottom_track_7 (
		.in({chanx_right_in[184], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_192_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_192_sram_inv[0:1]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_size2 mux_bottom_track_9 (
		.in({chanx_right_in[183], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_193_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_193_sram_inv[0:1]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size2 mux_bottom_track_11 (
		.in({chanx_right_in[182], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_194_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_194_sram_inv[0:1]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_size2 mux_bottom_track_13 (
		.in({chanx_right_in[181], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_195_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_195_sram_inv[0:1]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_size2 mux_bottom_track_15 (
		.in({chanx_right_in[180], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_196_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_196_sram_inv[0:1]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_size2 mux_bottom_track_17 (
		.in({chanx_right_in[179], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_197_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_197_sram_inv[0:1]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size2 mux_bottom_track_19 (
		.in({chanx_right_in[178], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_198_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_198_sram_inv[0:1]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_size2 mux_bottom_track_21 (
		.in({chanx_right_in[177], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_199_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_199_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_size2 mux_bottom_track_23 (
		.in({chanx_right_in[176], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_200_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_200_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_size2 mux_bottom_track_25 (
		.in({chanx_right_in[175], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_201_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_201_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size2 mux_bottom_track_27 (
		.in({chanx_right_in[174], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_202_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_202_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_size2 mux_bottom_track_29 (
		.in({chanx_right_in[173], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_203_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_203_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_size2 mux_bottom_track_31 (
		.in({chanx_right_in[172], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_204_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_204_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_size2 mux_bottom_track_33 (
		.in({chanx_right_in[171], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_205_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_205_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size2 mux_bottom_track_35 (
		.in({chanx_right_in[170], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_206_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_206_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_size2 mux_bottom_track_37 (
		.in({chanx_right_in[169], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_207_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_207_sram_inv[0:1]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_size2 mux_bottom_track_39 (
		.in({chanx_right_in[168], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_208_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_208_sram_inv[0:1]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_size2 mux_bottom_track_41 (
		.in({chanx_right_in[167], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_209_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_209_sram_inv[0:1]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size2 mux_bottom_track_43 (
		.in({chanx_right_in[166], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_210_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_210_sram_inv[0:1]),
		.out(chany_bottom_out[21]));

	mux_tree_tapbuf_size2 mux_bottom_track_45 (
		.in({chanx_right_in[165], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_211_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_211_sram_inv[0:1]),
		.out(chany_bottom_out[22]));

	mux_tree_tapbuf_size2 mux_bottom_track_47 (
		.in({chanx_right_in[164], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_212_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_212_sram_inv[0:1]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_size2 mux_bottom_track_49 (
		.in({chanx_right_in[163], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_213_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_213_sram_inv[0:1]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size2 mux_bottom_track_51 (
		.in({chanx_right_in[162], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_214_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_214_sram_inv[0:1]),
		.out(chany_bottom_out[25]));

	mux_tree_tapbuf_size2 mux_bottom_track_53 (
		.in({chanx_right_in[161], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_215_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_215_sram_inv[0:1]),
		.out(chany_bottom_out[26]));

	mux_tree_tapbuf_size2 mux_bottom_track_55 (
		.in({chanx_right_in[160], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_216_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_216_sram_inv[0:1]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_size2 mux_bottom_track_57 (
		.in({chanx_right_in[159], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_217_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_217_sram_inv[0:1]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size2 mux_bottom_track_59 (
		.in({chanx_right_in[158], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_218_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_218_sram_inv[0:1]),
		.out(chany_bottom_out[29]));

	mux_tree_tapbuf_size2 mux_bottom_track_61 (
		.in({chanx_right_in[157], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_219_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_219_sram_inv[0:1]),
		.out(chany_bottom_out[30]));

	mux_tree_tapbuf_size2 mux_bottom_track_63 (
		.in({chanx_right_in[156], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_220_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_220_sram_inv[0:1]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_size2 mux_bottom_track_65 (
		.in({chanx_right_in[155], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_221_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_221_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size2 mux_bottom_track_67 (
		.in({chanx_right_in[154], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_222_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_222_sram_inv[0:1]),
		.out(chany_bottom_out[33]));

	mux_tree_tapbuf_size2 mux_bottom_track_69 (
		.in({chanx_right_in[153], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_223_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_223_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	mux_tree_tapbuf_size2 mux_bottom_track_71 (
		.in({chanx_right_in[152], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_224_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_224_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	mux_tree_tapbuf_size2 mux_bottom_track_73 (
		.in({chanx_right_in[151], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_225_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_225_sram_inv[0:1]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size2 mux_bottom_track_75 (
		.in({chanx_right_in[150], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_226_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_226_sram_inv[0:1]),
		.out(chany_bottom_out[37]));

	mux_tree_tapbuf_size2 mux_bottom_track_77 (
		.in({chanx_right_in[149], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_227_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_227_sram_inv[0:1]),
		.out(chany_bottom_out[38]));

	mux_tree_tapbuf_size2 mux_bottom_track_79 (
		.in({chanx_right_in[148], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_228_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_228_sram_inv[0:1]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_size2 mux_bottom_track_81 (
		.in({chanx_right_in[147], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_229_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_229_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size2 mux_bottom_track_83 (
		.in({chanx_right_in[146], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_230_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_230_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	mux_tree_tapbuf_size2 mux_bottom_track_85 (
		.in({chanx_right_in[145], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_231_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_231_sram_inv[0:1]),
		.out(chany_bottom_out[42]));

	mux_tree_tapbuf_size2 mux_bottom_track_87 (
		.in({chanx_right_in[144], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_232_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_232_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	mux_tree_tapbuf_size2 mux_bottom_track_89 (
		.in({chanx_right_in[143], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_233_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_233_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size2 mux_bottom_track_91 (
		.in({chanx_right_in[142], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_234_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_234_sram_inv[0:1]),
		.out(chany_bottom_out[45]));

	mux_tree_tapbuf_size2 mux_bottom_track_93 (
		.in({chanx_right_in[141], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_235_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_235_sram_inv[0:1]),
		.out(chany_bottom_out[46]));

	mux_tree_tapbuf_size2 mux_bottom_track_95 (
		.in({chanx_right_in[140], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_236_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_236_sram_inv[0:1]),
		.out(chany_bottom_out[47]));

	mux_tree_tapbuf_size2 mux_bottom_track_97 (
		.in({chanx_right_in[139], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_237_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_237_sram_inv[0:1]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size2 mux_bottom_track_99 (
		.in({chanx_right_in[138], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_238_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_238_sram_inv[0:1]),
		.out(chany_bottom_out[49]));

	mux_tree_tapbuf_size2 mux_bottom_track_101 (
		.in({chanx_right_in[137], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_239_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_239_sram_inv[0:1]),
		.out(chany_bottom_out[50]));

	mux_tree_tapbuf_size2 mux_bottom_track_103 (
		.in({chanx_right_in[136], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_240_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_240_sram_inv[0:1]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_size2 mux_bottom_track_105 (
		.in({chanx_right_in[135], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_241_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_241_sram_inv[0:1]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size2 mux_bottom_track_107 (
		.in({chanx_right_in[134], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_242_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_242_sram_inv[0:1]),
		.out(chany_bottom_out[53]));

	mux_tree_tapbuf_size2 mux_bottom_track_109 (
		.in({chanx_right_in[133], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_243_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_243_sram_inv[0:1]),
		.out(chany_bottom_out[54]));

	mux_tree_tapbuf_size2 mux_bottom_track_111 (
		.in({chanx_right_in[132], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_244_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_244_sram_inv[0:1]),
		.out(chany_bottom_out[55]));

	mux_tree_tapbuf_size2 mux_bottom_track_113 (
		.in({chanx_right_in[131], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_245_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_245_sram_inv[0:1]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size2 mux_bottom_track_115 (
		.in({chanx_right_in[130], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_246_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_246_sram_inv[0:1]),
		.out(chany_bottom_out[57]));

	mux_tree_tapbuf_size2 mux_bottom_track_117 (
		.in({chanx_right_in[129], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_247_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_247_sram_inv[0:1]),
		.out(chany_bottom_out[58]));

	mux_tree_tapbuf_size2 mux_bottom_track_119 (
		.in({chanx_right_in[128], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_248_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_248_sram_inv[0:1]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_size2 mux_bottom_track_121 (
		.in({chanx_right_in[127], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_249_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_249_sram_inv[0:1]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size2 mux_bottom_track_123 (
		.in({chanx_right_in[126], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_250_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_250_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	mux_tree_tapbuf_size2 mux_bottom_track_125 (
		.in({chanx_right_in[125], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_251_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_251_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	mux_tree_tapbuf_size2 mux_bottom_track_127 (
		.in({chanx_right_in[124], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_252_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_252_sram_inv[0:1]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_size2 mux_bottom_track_129 (
		.in({chanx_right_in[123], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_253_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_253_sram_inv[0:1]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size2 mux_bottom_track_131 (
		.in({chanx_right_in[122], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_254_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_254_sram_inv[0:1]),
		.out(chany_bottom_out[65]));

	mux_tree_tapbuf_size2 mux_bottom_track_133 (
		.in({chanx_right_in[121], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_255_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_255_sram_inv[0:1]),
		.out(chany_bottom_out[66]));

	mux_tree_tapbuf_size2 mux_bottom_track_135 (
		.in({chanx_right_in[120], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_256_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_256_sram_inv[0:1]),
		.out(chany_bottom_out[67]));

	mux_tree_tapbuf_size2 mux_bottom_track_137 (
		.in({chanx_right_in[119], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_257_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_257_sram_inv[0:1]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size2 mux_bottom_track_139 (
		.in({chanx_right_in[118], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_258_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_258_sram_inv[0:1]),
		.out(chany_bottom_out[69]));

	mux_tree_tapbuf_size2 mux_bottom_track_141 (
		.in({chanx_right_in[117], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_259_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_259_sram_inv[0:1]),
		.out(chany_bottom_out[70]));

	mux_tree_tapbuf_size2 mux_bottom_track_143 (
		.in({chanx_right_in[116], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_260_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_260_sram_inv[0:1]),
		.out(chany_bottom_out[71]));

	mux_tree_tapbuf_size2 mux_bottom_track_145 (
		.in({chanx_right_in[115], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_261_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_261_sram_inv[0:1]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size2 mux_bottom_track_147 (
		.in({chanx_right_in[114], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_262_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_262_sram_inv[0:1]),
		.out(chany_bottom_out[73]));

	mux_tree_tapbuf_size2 mux_bottom_track_149 (
		.in({chanx_right_in[113], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_263_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_263_sram_inv[0:1]),
		.out(chany_bottom_out[74]));

	mux_tree_tapbuf_size2 mux_bottom_track_151 (
		.in({chanx_right_in[112], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_264_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_264_sram_inv[0:1]),
		.out(chany_bottom_out[75]));

	mux_tree_tapbuf_size2 mux_bottom_track_153 (
		.in({chanx_right_in[111], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_265_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_265_sram_inv[0:1]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size2 mux_bottom_track_155 (
		.in({chanx_right_in[110], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_266_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_266_sram_inv[0:1]),
		.out(chany_bottom_out[77]));

	mux_tree_tapbuf_size2 mux_bottom_track_157 (
		.in({chanx_right_in[109], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_267_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_267_sram_inv[0:1]),
		.out(chany_bottom_out[78]));

	mux_tree_tapbuf_size2 mux_bottom_track_159 (
		.in({chanx_right_in[108], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_268_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_268_sram_inv[0:1]),
		.out(chany_bottom_out[79]));

	mux_tree_tapbuf_size2 mux_bottom_track_161 (
		.in({chanx_right_in[107], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_269_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_269_sram_inv[0:1]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size2 mux_bottom_track_163 (
		.in({chanx_right_in[106], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_270_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_270_sram_inv[0:1]),
		.out(chany_bottom_out[81]));

	mux_tree_tapbuf_size2 mux_bottom_track_165 (
		.in({chanx_right_in[105], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_271_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_271_sram_inv[0:1]),
		.out(chany_bottom_out[82]));

	mux_tree_tapbuf_size2 mux_bottom_track_167 (
		.in({chanx_right_in[104], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_272_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_272_sram_inv[0:1]),
		.out(chany_bottom_out[83]));

	mux_tree_tapbuf_size2 mux_bottom_track_169 (
		.in({chanx_right_in[103], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_273_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_273_sram_inv[0:1]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size2 mux_bottom_track_171 (
		.in({chanx_right_in[102], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_274_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_274_sram_inv[0:1]),
		.out(chany_bottom_out[85]));

	mux_tree_tapbuf_size2 mux_bottom_track_173 (
		.in({chanx_right_in[101], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_275_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_275_sram_inv[0:1]),
		.out(chany_bottom_out[86]));

	mux_tree_tapbuf_size2 mux_bottom_track_175 (
		.in({chanx_right_in[100], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_276_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_276_sram_inv[0:1]),
		.out(chany_bottom_out[87]));

	mux_tree_tapbuf_size2 mux_bottom_track_177 (
		.in({chanx_right_in[99], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_277_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_277_sram_inv[0:1]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size2 mux_bottom_track_179 (
		.in({chanx_right_in[98], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_278_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_278_sram_inv[0:1]),
		.out(chany_bottom_out[89]));

	mux_tree_tapbuf_size2 mux_bottom_track_181 (
		.in({chanx_right_in[97], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_279_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_279_sram_inv[0:1]),
		.out(chany_bottom_out[90]));

	mux_tree_tapbuf_size2 mux_bottom_track_183 (
		.in({chanx_right_in[96], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_280_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_280_sram_inv[0:1]),
		.out(chany_bottom_out[91]));

	mux_tree_tapbuf_size2 mux_bottom_track_185 (
		.in({chanx_right_in[95], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_281_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_281_sram_inv[0:1]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size2 mux_bottom_track_187 (
		.in({chanx_right_in[94], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_282_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_282_sram_inv[0:1]),
		.out(chany_bottom_out[93]));

	mux_tree_tapbuf_size2 mux_bottom_track_189 (
		.in({chanx_right_in[93], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_283_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_283_sram_inv[0:1]),
		.out(chany_bottom_out[94]));

	mux_tree_tapbuf_size2 mux_bottom_track_191 (
		.in({chanx_right_in[92], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_284_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_284_sram_inv[0:1]),
		.out(chany_bottom_out[95]));

	mux_tree_tapbuf_size2 mux_bottom_track_193 (
		.in({chanx_right_in[91], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_285_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_285_sram_inv[0:1]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size2 mux_bottom_track_195 (
		.in({chanx_right_in[90], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_286_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_286_sram_inv[0:1]),
		.out(chany_bottom_out[97]));

	mux_tree_tapbuf_size2 mux_bottom_track_197 (
		.in({chanx_right_in[89], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_287_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_287_sram_inv[0:1]),
		.out(chany_bottom_out[98]));

	mux_tree_tapbuf_size2 mux_bottom_track_199 (
		.in({chanx_right_in[88], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_288_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_288_sram_inv[0:1]),
		.out(chany_bottom_out[99]));

	mux_tree_tapbuf_size2 mux_bottom_track_201 (
		.in({chanx_right_in[87], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_289_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_289_sram_inv[0:1]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size2 mux_bottom_track_203 (
		.in({chanx_right_in[86], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_290_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_290_sram_inv[0:1]),
		.out(chany_bottom_out[101]));

	mux_tree_tapbuf_size2 mux_bottom_track_205 (
		.in({chanx_right_in[85], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_291_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_291_sram_inv[0:1]),
		.out(chany_bottom_out[102]));

	mux_tree_tapbuf_size2 mux_bottom_track_207 (
		.in({chanx_right_in[84], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_292_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_292_sram_inv[0:1]),
		.out(chany_bottom_out[103]));

	mux_tree_tapbuf_size2 mux_bottom_track_209 (
		.in({chanx_right_in[83], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_293_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_293_sram_inv[0:1]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size2 mux_bottom_track_211 (
		.in({chanx_right_in[82], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_294_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_294_sram_inv[0:1]),
		.out(chany_bottom_out[105]));

	mux_tree_tapbuf_size2 mux_bottom_track_213 (
		.in({chanx_right_in[81], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_295_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_295_sram_inv[0:1]),
		.out(chany_bottom_out[106]));

	mux_tree_tapbuf_size2 mux_bottom_track_215 (
		.in({chanx_right_in[80], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_296_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_296_sram_inv[0:1]),
		.out(chany_bottom_out[107]));

	mux_tree_tapbuf_size2 mux_bottom_track_217 (
		.in({chanx_right_in[79], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_297_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_297_sram_inv[0:1]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size2 mux_bottom_track_219 (
		.in({chanx_right_in[78], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_298_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_298_sram_inv[0:1]),
		.out(chany_bottom_out[109]));

	mux_tree_tapbuf_size2 mux_bottom_track_221 (
		.in({chanx_right_in[77], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_299_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_299_sram_inv[0:1]),
		.out(chany_bottom_out[110]));

	mux_tree_tapbuf_size2 mux_bottom_track_223 (
		.in({chanx_right_in[76], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_300_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_300_sram_inv[0:1]),
		.out(chany_bottom_out[111]));

	mux_tree_tapbuf_size2 mux_bottom_track_225 (
		.in({chanx_right_in[75], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_301_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_301_sram_inv[0:1]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size2 mux_bottom_track_227 (
		.in({chanx_right_in[74], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_302_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_302_sram_inv[0:1]),
		.out(chany_bottom_out[113]));

	mux_tree_tapbuf_size2 mux_bottom_track_229 (
		.in({chanx_right_in[73], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_303_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_303_sram_inv[0:1]),
		.out(chany_bottom_out[114]));

	mux_tree_tapbuf_size2 mux_bottom_track_231 (
		.in({chanx_right_in[72], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_304_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_304_sram_inv[0:1]),
		.out(chany_bottom_out[115]));

	mux_tree_tapbuf_size2 mux_bottom_track_233 (
		.in({chanx_right_in[71], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_305_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_305_sram_inv[0:1]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size2 mux_bottom_track_235 (
		.in({chanx_right_in[70], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_306_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_306_sram_inv[0:1]),
		.out(chany_bottom_out[117]));

	mux_tree_tapbuf_size2 mux_bottom_track_237 (
		.in({chanx_right_in[69], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_307_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_307_sram_inv[0:1]),
		.out(chany_bottom_out[118]));

	mux_tree_tapbuf_size2 mux_bottom_track_239 (
		.in({chanx_right_in[68], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_308_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_308_sram_inv[0:1]),
		.out(chany_bottom_out[119]));

	mux_tree_tapbuf_size2 mux_bottom_track_241 (
		.in({chanx_right_in[67], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_309_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_309_sram_inv[0:1]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size2 mux_bottom_track_243 (
		.in({chanx_right_in[66], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_310_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_310_sram_inv[0:1]),
		.out(chany_bottom_out[121]));

	mux_tree_tapbuf_size2 mux_bottom_track_245 (
		.in({chanx_right_in[65], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_311_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_311_sram_inv[0:1]),
		.out(chany_bottom_out[122]));

	mux_tree_tapbuf_size2 mux_bottom_track_247 (
		.in({chanx_right_in[64], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_312_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_312_sram_inv[0:1]),
		.out(chany_bottom_out[123]));

	mux_tree_tapbuf_size2 mux_bottom_track_249 (
		.in({chanx_right_in[63], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_313_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_313_sram_inv[0:1]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size2 mux_bottom_track_251 (
		.in({chanx_right_in[62], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_314_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_314_sram_inv[0:1]),
		.out(chany_bottom_out[125]));

	mux_tree_tapbuf_size2 mux_bottom_track_253 (
		.in({chanx_right_in[61], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_315_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_315_sram_inv[0:1]),
		.out(chany_bottom_out[126]));

	mux_tree_tapbuf_size2 mux_bottom_track_255 (
		.in({chanx_right_in[60], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_316_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_316_sram_inv[0:1]),
		.out(chany_bottom_out[127]));

	mux_tree_tapbuf_size2 mux_bottom_track_257 (
		.in({chanx_right_in[59], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_317_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_317_sram_inv[0:1]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size2 mux_bottom_track_259 (
		.in({chanx_right_in[58], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_318_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_318_sram_inv[0:1]),
		.out(chany_bottom_out[129]));

	mux_tree_tapbuf_size2 mux_bottom_track_261 (
		.in({chanx_right_in[57], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_319_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_319_sram_inv[0:1]),
		.out(chany_bottom_out[130]));

	mux_tree_tapbuf_size2 mux_bottom_track_263 (
		.in({chanx_right_in[56], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_320_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_320_sram_inv[0:1]),
		.out(chany_bottom_out[131]));

	mux_tree_tapbuf_size2 mux_bottom_track_265 (
		.in({chanx_right_in[55], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_321_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_321_sram_inv[0:1]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size2 mux_bottom_track_267 (
		.in({chanx_right_in[54], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_322_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_322_sram_inv[0:1]),
		.out(chany_bottom_out[133]));

	mux_tree_tapbuf_size2 mux_bottom_track_269 (
		.in({chanx_right_in[53], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_323_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_323_sram_inv[0:1]),
		.out(chany_bottom_out[134]));

	mux_tree_tapbuf_size2 mux_bottom_track_271 (
		.in({chanx_right_in[52], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_324_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_324_sram_inv[0:1]),
		.out(chany_bottom_out[135]));

	mux_tree_tapbuf_size2 mux_bottom_track_273 (
		.in({chanx_right_in[51], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_325_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_325_sram_inv[0:1]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size2 mux_bottom_track_275 (
		.in({chanx_right_in[50], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_326_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_326_sram_inv[0:1]),
		.out(chany_bottom_out[137]));

	mux_tree_tapbuf_size2 mux_bottom_track_277 (
		.in({chanx_right_in[49], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_327_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_327_sram_inv[0:1]),
		.out(chany_bottom_out[138]));

	mux_tree_tapbuf_size2 mux_bottom_track_279 (
		.in({chanx_right_in[48], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_328_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_328_sram_inv[0:1]),
		.out(chany_bottom_out[139]));

	mux_tree_tapbuf_size2 mux_bottom_track_281 (
		.in({chanx_right_in[47], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_329_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_329_sram_inv[0:1]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size2 mux_bottom_track_283 (
		.in({chanx_right_in[46], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_330_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_330_sram_inv[0:1]),
		.out(chany_bottom_out[141]));

	mux_tree_tapbuf_size2 mux_bottom_track_285 (
		.in({chanx_right_in[45], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_331_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_331_sram_inv[0:1]),
		.out(chany_bottom_out[142]));

	mux_tree_tapbuf_size2 mux_bottom_track_287 (
		.in({chanx_right_in[44], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_332_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_332_sram_inv[0:1]),
		.out(chany_bottom_out[143]));

	mux_tree_tapbuf_size2 mux_bottom_track_289 (
		.in({chanx_right_in[43], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_333_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_333_sram_inv[0:1]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size2 mux_bottom_track_291 (
		.in({chanx_right_in[42], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_334_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_334_sram_inv[0:1]),
		.out(chany_bottom_out[145]));

	mux_tree_tapbuf_size2 mux_bottom_track_293 (
		.in({chanx_right_in[41], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_335_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_335_sram_inv[0:1]),
		.out(chany_bottom_out[146]));

	mux_tree_tapbuf_size2 mux_bottom_track_295 (
		.in({chanx_right_in[40], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_336_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_336_sram_inv[0:1]),
		.out(chany_bottom_out[147]));

	mux_tree_tapbuf_size2 mux_bottom_track_297 (
		.in({chanx_right_in[39], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_337_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_337_sram_inv[0:1]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size2 mux_bottom_track_299 (
		.in({chanx_right_in[38], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_338_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_338_sram_inv[0:1]),
		.out(chany_bottom_out[149]));

	mux_tree_tapbuf_size2 mux_bottom_track_301 (
		.in({chanx_right_in[37], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_339_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_339_sram_inv[0:1]),
		.out(chany_bottom_out[150]));

	mux_tree_tapbuf_size2 mux_bottom_track_303 (
		.in({chanx_right_in[36], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_340_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_340_sram_inv[0:1]),
		.out(chany_bottom_out[151]));

	mux_tree_tapbuf_size2 mux_bottom_track_305 (
		.in({chanx_right_in[35], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_341_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_341_sram_inv[0:1]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size2 mux_bottom_track_307 (
		.in({chanx_right_in[34], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_342_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_342_sram_inv[0:1]),
		.out(chany_bottom_out[153]));

	mux_tree_tapbuf_size2 mux_bottom_track_309 (
		.in({chanx_right_in[33], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_343_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_343_sram_inv[0:1]),
		.out(chany_bottom_out[154]));

	mux_tree_tapbuf_size2 mux_bottom_track_311 (
		.in({chanx_right_in[32], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_344_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_344_sram_inv[0:1]),
		.out(chany_bottom_out[155]));

	mux_tree_tapbuf_size2 mux_bottom_track_313 (
		.in({chanx_right_in[31], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_345_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_345_sram_inv[0:1]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size2 mux_bottom_track_315 (
		.in({chanx_right_in[30], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_346_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_346_sram_inv[0:1]),
		.out(chany_bottom_out[157]));

	mux_tree_tapbuf_size2 mux_bottom_track_317 (
		.in({chanx_right_in[29], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_347_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_347_sram_inv[0:1]),
		.out(chany_bottom_out[158]));

	mux_tree_tapbuf_size2 mux_bottom_track_319 (
		.in({chanx_right_in[28], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_348_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_348_sram_inv[0:1]),
		.out(chany_bottom_out[159]));

	mux_tree_tapbuf_size2 mux_bottom_track_321 (
		.in({chanx_right_in[27], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_349_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_349_sram_inv[0:1]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size2 mux_bottom_track_323 (
		.in({chanx_right_in[26], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_350_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_350_sram_inv[0:1]),
		.out(chany_bottom_out[161]));

	mux_tree_tapbuf_size2 mux_bottom_track_325 (
		.in({chanx_right_in[25], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_351_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_351_sram_inv[0:1]),
		.out(chany_bottom_out[162]));

	mux_tree_tapbuf_size2 mux_bottom_track_327 (
		.in({chanx_right_in[24], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_352_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_352_sram_inv[0:1]),
		.out(chany_bottom_out[163]));

	mux_tree_tapbuf_size2 mux_bottom_track_329 (
		.in({chanx_right_in[23], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_353_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_353_sram_inv[0:1]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size2 mux_bottom_track_331 (
		.in({chanx_right_in[22], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_354_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_354_sram_inv[0:1]),
		.out(chany_bottom_out[165]));

	mux_tree_tapbuf_size2 mux_bottom_track_333 (
		.in({chanx_right_in[21], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_355_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_355_sram_inv[0:1]),
		.out(chany_bottom_out[166]));

	mux_tree_tapbuf_size2 mux_bottom_track_335 (
		.in({chanx_right_in[20], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_356_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_356_sram_inv[0:1]),
		.out(chany_bottom_out[167]));

	mux_tree_tapbuf_size2 mux_bottom_track_337 (
		.in({chanx_right_in[19], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_357_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_357_sram_inv[0:1]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size2 mux_bottom_track_339 (
		.in({chanx_right_in[18], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_358_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_358_sram_inv[0:1]),
		.out(chany_bottom_out[169]));

	mux_tree_tapbuf_size2 mux_bottom_track_341 (
		.in({chanx_right_in[17], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_359_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_359_sram_inv[0:1]),
		.out(chany_bottom_out[170]));

	mux_tree_tapbuf_size2 mux_bottom_track_343 (
		.in({chanx_right_in[16], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_360_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_360_sram_inv[0:1]),
		.out(chany_bottom_out[171]));

	mux_tree_tapbuf_size2 mux_bottom_track_345 (
		.in({chanx_right_in[15], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_361_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_361_sram_inv[0:1]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size2 mux_bottom_track_347 (
		.in({chanx_right_in[14], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_362_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_362_sram_inv[0:1]),
		.out(chany_bottom_out[173]));

	mux_tree_tapbuf_size2 mux_bottom_track_349 (
		.in({chanx_right_in[13], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_363_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_363_sram_inv[0:1]),
		.out(chany_bottom_out[174]));

	mux_tree_tapbuf_size2 mux_bottom_track_351 (
		.in({chanx_right_in[12], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_364_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_364_sram_inv[0:1]),
		.out(chany_bottom_out[175]));

	mux_tree_tapbuf_size2 mux_bottom_track_353 (
		.in({chanx_right_in[11], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_365_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_365_sram_inv[0:1]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size2 mux_bottom_track_355 (
		.in({chanx_right_in[10], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_366_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_366_sram_inv[0:1]),
		.out(chany_bottom_out[177]));

	mux_tree_tapbuf_size2 mux_bottom_track_357 (
		.in({chanx_right_in[9], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_367_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_367_sram_inv[0:1]),
		.out(chany_bottom_out[178]));

	mux_tree_tapbuf_size2 mux_bottom_track_359 (
		.in({chanx_right_in[8], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_368_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_368_sram_inv[0:1]),
		.out(chany_bottom_out[179]));

	mux_tree_tapbuf_size2 mux_bottom_track_361 (
		.in({chanx_right_in[7], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size2_369_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_369_sram_inv[0:1]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size2 mux_bottom_track_363 (
		.in({chanx_right_in[6], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_370_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_370_sram_inv[0:1]),
		.out(chany_bottom_out[181]));

	mux_tree_tapbuf_size2 mux_bottom_track_365 (
		.in({chanx_right_in[5], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_371_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_371_sram_inv[0:1]),
		.out(chany_bottom_out[182]));

	mux_tree_tapbuf_size2 mux_bottom_track_367 (
		.in({chanx_right_in[4], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_372_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_372_sram_inv[0:1]),
		.out(chany_bottom_out[183]));

	mux_tree_tapbuf_size2 mux_bottom_track_369 (
		.in({chanx_right_in[3], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_373_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_373_sram_inv[0:1]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size2 mux_bottom_track_371 (
		.in({chanx_right_in[2], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_374_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_374_sram_inv[0:1]),
		.out(chany_bottom_out[185]));

	mux_tree_tapbuf_size2 mux_bottom_track_373 (
		.in({chanx_right_in[1], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_375_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_375_sram_inv[0:1]),
		.out(chany_bottom_out[186]));

	mux_tree_tapbuf_size2 mux_bottom_track_375 (
		.in({chanx_right_in[0], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_376_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_376_sram_inv[0:1]),
		.out(chany_bottom_out[187]));

	mux_tree_tapbuf_size2 mux_bottom_track_377 (
		.in({chanx_right_in[188], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_377_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_377_sram_inv[0:1]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size2_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_27_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_28_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_29_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_30_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_31_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_32_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_33_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_34_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_35_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_36_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_37_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_38_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_39_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_40_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_41_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_42_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_43_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_44_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_45_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_46_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_47_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_48_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_49_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_50_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_51_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_52_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_53_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_54_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_55_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_56_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_57_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_58_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_59_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_60_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_61_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_62_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_63_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_64_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_65_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_66_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_67_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_68_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_69_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_70_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_71_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_72_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_73_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_74_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_75_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_76_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_77_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_78_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_79_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_80_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_81_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_82_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_83_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_84_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_85_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_86_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_87_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_88_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_89_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_90_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_91_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_92_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_93_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_94_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_95_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_96_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_97_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_98_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_99_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_100_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_101_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_102_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_103_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_104_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_105_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_212 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_106_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_214 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_107_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_108_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_218 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_109_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_220 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_110_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_222 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_111_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_112_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_226 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_113_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_228 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_114_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_230 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_115_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_116_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_234 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_117_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_236 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_118_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_238 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_119_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_120_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_120_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_242 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_121_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_121_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_244 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_122_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_122_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_246 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_123_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_123_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_124_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_124_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_250 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_125_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_125_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_252 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_126_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_126_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_254 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_127_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_127_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_128_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_128_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_258 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_129_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_129_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_260 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_130_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_130_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_262 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_131_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_131_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_132_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_132_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_266 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_133_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_133_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_268 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_134_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_134_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_270 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_135_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_135_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_136_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_136_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_136_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_274 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_136_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_137_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_137_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_137_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_276 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_137_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_138_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_138_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_138_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_278 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_138_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_139_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_139_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_139_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_139_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_140_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_140_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_140_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_282 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_140_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_141_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_141_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_141_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_284 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_141_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_142_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_142_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_142_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_286 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_142_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_143_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_143_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_143_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_143_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_144_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_144_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_144_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_290 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_144_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_145_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_145_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_145_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_292 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_145_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_146_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_146_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_146_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_294 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_146_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_147_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_147_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_147_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_147_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_148_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_148_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_148_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_298 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_148_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_149_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_149_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_149_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_300 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_149_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_150_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_150_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_150_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_302 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_150_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_151_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_151_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_151_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_151_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_152_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_152_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_152_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_306 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_152_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_153_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_153_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_153_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_308 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_153_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_154_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_154_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_154_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_310 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_154_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_155_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_155_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_155_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_155_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_156_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_156_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_156_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_314 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_156_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_157_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_157_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_157_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_316 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_157_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_158_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_158_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_158_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_318 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_158_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_159_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_159_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_159_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_159_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_160_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_160_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_160_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_322 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_160_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_161_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_161_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_161_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_324 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_161_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_162_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_162_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_162_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_326 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_162_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_163_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_163_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_163_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_163_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_164_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_164_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_164_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_330 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_164_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_165_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_165_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_165_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_332 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_165_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_166_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_166_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_166_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_334 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_166_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_167_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_167_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_167_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_167_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_168_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_168_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_168_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_338 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_168_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_169_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_169_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_169_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_340 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_169_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_170_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_170_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_170_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_342 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_170_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_171_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_171_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_171_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_171_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_172_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_172_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_172_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_346 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_172_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_173_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_173_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_173_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_348 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_173_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_174_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_174_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_174_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_350 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_174_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_175_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_175_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_175_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_175_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_176_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_176_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_176_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_354 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_176_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_177_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_177_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_177_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_356 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_177_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_178_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_178_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_178_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_358 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_178_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_179_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_179_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_179_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_179_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_180_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_180_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_180_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_362 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_180_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_181_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_181_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_181_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_364 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_181_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_182_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_182_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_182_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_366 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_182_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_183_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_183_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_183_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_183_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_184_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_184_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_184_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_370 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_184_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_185_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_185_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_185_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_372 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_185_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_186_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_186_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_186_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_374 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_186_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_187_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_187_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_187_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_187_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_188_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_188_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_188_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_188_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_189_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_189_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_189_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_189_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_190_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_190_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_190_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_190_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_191_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_191_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_191_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_191_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_192_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_192_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_192_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_192_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_193_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_193_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_193_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_193_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_194_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_194_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_194_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_194_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_195_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_195_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_195_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_195_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_196_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_196_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_196_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_196_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_197_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_197_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_197_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_197_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_198_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_198_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_198_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_198_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_199_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_199_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_199_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_199_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_200_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_200_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_200_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_200_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_201_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_201_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_201_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_201_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_202_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_202_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_202_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_202_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_203_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_203_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_203_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_203_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_204_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_204_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_204_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_204_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_205_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_205_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_205_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_205_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_206_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_206_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_206_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_206_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_207_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_207_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_207_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_207_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_208_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_208_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_208_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_208_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_209_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_209_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_209_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_209_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_210_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_210_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_210_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_210_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_211_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_211_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_211_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_211_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_212_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_212_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_212_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_212_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_213_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_213_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_213_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_213_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_214_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_214_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_214_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_214_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_215_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_215_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_215_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_215_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_216_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_216_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_216_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_216_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_217_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_217_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_217_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_217_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_218_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_218_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_218_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_218_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_219_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_219_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_219_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_219_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_220_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_220_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_220_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_220_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_221_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_221_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_221_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_221_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_222_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_222_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_222_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_222_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_223_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_223_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_223_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_223_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_224_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_224_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_224_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_224_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_225_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_225_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_225_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_225_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_226_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_226_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_226_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_226_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_227_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_227_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_227_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_227_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_228_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_228_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_228_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_228_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_229_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_229_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_229_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_229_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_230_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_230_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_230_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_230_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_231_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_231_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_231_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_231_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_232_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_232_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_232_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_232_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_233_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_233_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_233_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_233_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_234_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_234_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_234_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_234_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_235_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_235_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_235_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_235_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_236_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_236_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_236_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_236_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_237_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_237_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_237_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_237_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_238_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_238_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_238_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_238_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_239_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_239_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_239_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_239_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_240_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_240_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_240_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_240_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_241_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_241_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_241_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_241_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_242_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_242_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_242_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_242_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_243_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_243_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_243_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_243_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_244_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_244_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_244_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_244_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_245_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_245_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_245_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_245_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_246_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_246_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_246_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_246_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_247_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_247_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_247_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_247_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_248_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_248_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_248_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_248_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_249_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_249_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_249_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_249_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_250_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_250_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_250_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_250_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_251_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_251_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_251_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_251_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_252_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_252_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_252_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_252_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_253_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_253_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_253_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_253_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_254_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_254_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_254_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_254_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_255_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_255_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_255_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_255_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_256_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_256_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_256_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_256_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_257_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_257_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_257_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_257_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_258_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_258_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_258_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_258_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_259_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_259_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_259_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_259_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_260_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_260_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_260_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_260_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_261_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_261_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_261_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_147 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_261_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_262_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_262_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_262_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_149 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_262_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_263_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_263_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_263_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_151 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_263_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_264_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_264_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_264_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_264_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_265_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_265_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_265_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_155 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_265_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_266_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_266_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_266_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_157 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_266_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_267_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_267_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_267_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_159 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_267_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_268_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_268_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_268_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_268_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_269_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_269_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_269_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_163 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_269_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_270_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_270_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_270_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_165 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_270_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_271_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_271_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_271_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_167 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_271_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_272_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_272_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_272_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_272_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_273_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_273_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_273_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_171 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_273_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_274_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_274_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_274_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_173 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_274_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_275_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_275_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_275_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_175 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_275_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_276_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_276_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_276_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_276_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_277_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_277_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_277_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_179 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_277_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_278_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_278_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_278_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_181 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_278_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_279_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_279_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_279_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_183 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_279_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_280_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_280_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_280_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_280_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_281_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_281_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_281_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_187 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_281_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_282_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_282_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_282_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_189 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_282_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_283_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_283_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_283_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_191 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_283_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_284_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_284_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_284_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_284_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_285_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_285_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_285_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_195 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_285_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_286_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_286_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_286_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_197 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_286_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_287_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_287_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_287_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_199 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_287_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_288_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_288_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_288_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_288_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_289_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_289_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_289_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_203 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_289_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_290_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_290_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_290_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_205 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_290_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_291_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_291_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_291_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_207 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_291_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_292_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_292_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_292_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_292_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_293_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_293_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_293_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_211 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_293_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_294_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_294_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_294_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_213 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_294_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_295_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_295_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_295_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_215 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_295_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_296_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_296_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_296_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_296_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_297_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_297_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_297_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_219 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_297_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_298_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_298_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_298_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_221 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_298_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_299_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_299_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_299_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_223 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_299_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_300_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_300_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_300_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_300_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_301_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_301_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_301_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_227 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_301_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_302_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_302_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_302_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_229 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_302_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_303_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_303_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_303_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_231 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_303_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_304_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_304_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_304_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_304_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_305_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_305_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_305_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_235 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_305_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_306_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_306_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_306_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_237 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_306_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_307_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_307_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_307_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_239 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_307_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_308_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_308_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_308_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_308_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_309_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_309_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_309_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_243 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_309_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_310_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_310_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_310_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_245 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_310_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_311_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_311_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_311_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_247 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_311_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_312_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_312_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_312_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_312_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_313_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_313_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_313_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_251 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_313_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_314_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_314_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_314_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_253 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_314_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_315_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_315_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_315_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_255 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_315_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_316_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_316_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_316_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_316_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_317_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_317_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_317_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_259 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_317_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_318_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_318_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_318_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_261 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_318_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_319_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_319_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_319_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_263 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_319_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_320_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_320_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_320_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_320_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_321_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_321_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_321_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_267 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_321_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_322_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_322_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_322_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_269 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_322_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_323_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_323_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_323_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_271 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_323_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_324_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_324_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_324_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_324_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_325_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_325_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_325_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_275 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_325_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_326_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_326_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_326_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_277 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_326_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_327_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_327_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_327_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_279 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_327_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_328_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_328_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_328_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_328_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_329_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_329_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_329_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_283 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_329_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_330_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_330_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_330_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_285 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_330_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_331_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_331_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_331_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_287 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_331_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_332_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_332_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_332_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_332_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_333_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_333_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_333_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_291 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_333_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_334_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_334_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_334_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_293 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_334_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_335_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_335_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_335_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_295 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_335_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_336_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_336_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_336_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_336_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_337_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_337_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_337_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_299 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_337_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_338_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_338_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_338_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_301 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_338_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_339_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_339_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_339_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_303 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_339_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_340_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_340_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_340_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_340_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_341_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_341_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_341_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_307 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_341_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_342_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_342_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_342_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_309 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_342_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_343_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_343_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_343_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_311 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_343_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_344_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_344_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_344_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_344_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_345_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_345_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_345_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_315 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_345_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_346_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_346_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_346_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_317 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_346_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_347_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_347_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_347_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_319 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_347_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_348_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_348_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_348_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_348_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_349_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_349_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_349_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_323 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_349_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_350_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_350_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_350_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_325 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_350_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_351_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_351_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_351_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_327 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_351_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_352_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_352_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_352_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_352_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_353_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_353_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_353_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_331 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_353_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_354_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_354_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_354_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_333 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_354_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_355_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_355_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_355_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_335 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_355_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_356_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_356_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_356_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_356_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_357_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_357_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_357_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_339 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_357_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_358_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_358_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_358_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_341 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_358_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_359_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_359_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_359_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_343 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_359_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_360_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_360_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_360_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_360_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_361_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_361_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_361_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_347 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_361_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_362_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_362_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_362_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_349 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_362_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_363_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_363_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_363_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_351 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_363_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_364_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_364_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_364_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_364_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_365_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_365_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_365_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_355 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_365_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_366_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_366_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_366_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_357 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_366_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_367_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_367_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_367_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_359 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_367_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_368_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_368_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_368_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_368_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_369_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_369_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_369_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_363 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_369_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_370_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_370_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_370_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_365 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_370_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_371_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_371_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_371_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_367 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_371_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_372_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_372_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_372_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_372_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_373_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_373_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_373_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_371 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_373_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_374_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_374_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_374_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_373 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_374_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_375_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_375_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_375_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_375 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_375_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_376_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_376_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_376_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_376_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_377_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_377_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_0__6_ -----

//----- Default net type -----
`default_nettype wire



