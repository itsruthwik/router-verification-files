//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: router_tb
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jun 28 12:51:29 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

module router_tb_top_formal_verification (
input [0:0] clk,
input [0:0] reset,
input [0:0] router_address_5_,
input [0:0] router_address_4_,
input [0:0] router_address_3_,
input [0:0] router_address_2_,
input [0:0] router_address_1_,
input [0:0] router_address_0_,
output [0:0] rtr_error);

// ----- Local wires for FPGA fabric -----
wire [0:159] gfpga_pad_GPIO_PAD_fm;
wire [0:0] ccff_head_fm;
wire [0:0] ccff_tail_fm;
wire [0:0] prog_clk_fm;
wire [0:0] set_fm;
wire [0:0] reset_fm;
wire [0:0] clk_fm;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		prog_clk_fm[0],
		set_fm[0],
		reset_fm[0],
		clk_fm[0],
		gfpga_pad_GPIO_PAD_fm[0:159],
		ccff_head_fm[0],
		ccff_tail_fm[0]);

// ----- Begin Connect Global ports of FPGA top module -----
	assign set_fm[0] = 1'b0;
	assign reset_fm[0] = 1'b0;
	assign clk_fm[0] = clk[0];
	assign prog_clk_fm[0] = 1'b0;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input clk is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[127] -----
	assign gfpga_pad_GPIO_PAD_fm[127] = clk[0];

// ----- Blif Benchmark input reset is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[121] -----
	assign gfpga_pad_GPIO_PAD_fm[121] = reset[0];

// ----- Blif Benchmark input router_address_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[124] -----
	assign gfpga_pad_GPIO_PAD_fm[124] = router_address_5_[0];

// ----- Blif Benchmark input router_address_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[126] -----
	assign gfpga_pad_GPIO_PAD_fm[126] = router_address_4_[0];

// ----- Blif Benchmark input router_address_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[122] -----
	assign gfpga_pad_GPIO_PAD_fm[122] = router_address_3_[0];

// ----- Blif Benchmark input router_address_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[120] -----
	assign gfpga_pad_GPIO_PAD_fm[120] = router_address_2_[0];

// ----- Blif Benchmark input router_address_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[123] -----
	assign gfpga_pad_GPIO_PAD_fm[123] = router_address_1_[0];

// ----- Blif Benchmark input router_address_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[128] -----
	assign gfpga_pad_GPIO_PAD_fm[128] = router_address_0_[0];

// ----- Blif Benchmark output rtr_error is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[138] -----
	assign rtr_error[0] = gfpga_pad_GPIO_PAD_fm[138];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD_fm[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[2] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[3] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[4] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[6] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[7] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[11] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[12] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[14] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[26] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[31] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[32] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[33] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[34] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[35] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[36] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[37] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[38] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[39] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[40] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[41] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[42] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[43] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[44] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[45] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[46] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[47] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[48] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[49] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[50] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[51] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[52] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[53] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[54] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[55] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[56] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[57] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[58] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[59] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[60] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[61] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[62] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[63] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[64] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[65] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[66] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[67] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[68] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[69] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[70] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[71] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[72] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[73] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[74] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[75] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[76] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[77] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[78] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[79] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[80] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[81] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[82] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[83] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[84] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[85] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[86] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[87] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[88] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[89] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[90] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[91] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[92] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[93] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[94] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[95] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[96] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[97] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[98] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[99] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[100] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[101] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[102] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[103] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[104] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[105] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[106] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[107] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[108] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[109] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[110] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[111] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[112] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[113] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[114] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[115] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[116] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[117] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[118] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[119] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[125] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[129] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[130] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[131] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[132] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[133] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[134] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[135] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[136] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[137] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[139] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[140] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[141] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[142] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[143] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[144] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[145] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[146] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[147] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[148] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[149] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[150] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[151] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[152] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[153] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[154] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[155] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[156] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[157] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[158] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[159] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
// ----- Begin assign bitstream to configuration memories -----
initial begin
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b0000000011111111;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b1111111100000000;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b0101010110101010;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b1010101001010101;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b0101111110100000;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b1010000001011111;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b0110101010101010;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b1001010101010101;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b0011001111001100;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b1100110000110011;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b1000000000000000;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b0111111111111111;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b0011110011110000;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b1100001100001111;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b1110111011101110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b0001000100010001;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_210.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_210.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_212.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_212.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_216.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_216.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_218.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_218.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_222.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_222.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_224.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_224.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_226.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_226.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_228.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_228.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_234.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_234.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_236.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_236.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_240.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_240.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_244.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_244.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_248.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_248.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_252.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_252.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_256.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_256.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_258.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_258.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_260.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_260.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_266.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_266.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_270.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_270.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_272.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_272.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_274.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_274.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_276.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_276.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_280.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_280.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_284.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_284.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_288.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_288.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_290.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_290.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_296.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_296.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_298.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_298.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_300.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_300.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_306.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_306.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_308.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_308.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_312.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_312.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_314.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_314.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_316.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_316.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_320.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_320.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_324.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_324.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_328.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_328.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_330.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_330.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_332.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_332.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_336.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_336.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_338.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_338.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_342.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_342.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_344.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_344.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_346.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_346.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_348.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_348.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_352.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_352.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_354.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_354.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_356.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_356.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_360.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_360.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_362.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_362.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_364.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_364.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_368.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_368.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_370.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_370.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_372.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_372.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_376.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_376.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_378.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_378.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_380.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_380.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_384.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_384.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_76.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_76.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_84.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_84.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_92.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_92.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_108.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_108.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_116.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_116.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_124.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_124.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_132.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_132.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_140.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_140.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_148.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_148.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_156.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_156.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_172.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_172.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_180.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_180.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_186.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_186.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_188.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_188.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_204.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_204.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_210.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_210.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_212.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_212.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_214.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_214.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_216.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_216.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_218.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_218.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_222.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_222.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_224.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_224.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_226.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_226.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_228.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_228.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_232.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_232.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_234.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_234.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_236.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_236.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_240.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_240.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_244.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_244.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_248.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_248.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_250.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_250.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_252.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_252.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_256.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_256.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_258.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_258.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_260.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_260.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_266.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_266.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_268.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_268.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_270.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_270.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_272.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_272.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_274.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_274.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_276.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_276.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_280.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_280.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_284.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_284.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_286.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_286.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_288.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_288.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_290.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_290.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_296.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_296.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_298.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_298.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_300.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_300.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_304.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_304.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_306.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_306.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_308.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_308.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_312.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_312.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_314.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_314.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_316.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_316.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_320.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_320.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_322.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_322.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_324.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_324.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_328.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_328.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_330.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_330.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_332.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_332.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_336.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_336.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_338.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_338.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_340.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_340.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_342.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_342.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_344.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_344.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_346.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_346.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_348.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_348.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_352.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_352.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_354.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_354.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_356.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_356.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_358.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_358.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_360.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_360.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_362.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_362.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_364.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_364.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_368.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_368.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_370.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_370.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_372.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_372.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_376.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_376.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_378.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_378.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_380.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_380.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_384.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_384.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__1_.mem_top_track_72.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_0__1_.mem_top_track_72.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_0__1_.mem_top_track_80.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__1_.mem_top_track_80.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__1_.mem_top_track_88.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__1_.mem_top_track_88.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__1_.mem_top_track_96.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__1_.mem_top_track_96.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__1_.mem_top_track_104.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__1_.mem_top_track_104.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__1_.mem_top_track_112.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__1_.mem_top_track_112.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__1_.mem_top_track_120.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__1_.mem_top_track_120.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__1_.mem_top_track_128.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_0__1_.mem_top_track_128.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_0__1_.mem_top_track_136.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_0__1_.mem_top_track_136.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_0__1_.mem_top_track_144.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__1_.mem_top_track_144.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__1_.mem_top_track_152.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__1_.mem_top_track_152.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__1_.mem_top_track_160.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__1_.mem_top_track_160.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__1_.mem_top_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_176.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__1_.mem_top_track_176.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__1_.mem_top_track_184.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_0__1_.mem_top_track_184.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_0__1_.mem_top_track_192.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__1_.mem_top_track_192.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__1_.mem_top_track_200.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__1_.mem_top_track_200.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__1_.mem_top_track_208.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_208.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_216.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__1_.mem_top_track_216.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__1_.mem_top_track_224.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_0__1_.mem_top_track_224.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_0__1_.mem_top_track_232.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__1_.mem_top_track_232.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__1_.mem_top_track_240.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_0__1_.mem_top_track_240.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_0__1_.mem_top_track_248.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_0__1_.mem_top_track_248.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_0__1_.mem_top_track_256.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__1_.mem_top_track_256.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__1_.mem_top_track_264.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__1_.mem_top_track_264.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__1_.mem_top_track_272.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__1_.mem_top_track_272.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__1_.mem_top_track_280.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__1_.mem_top_track_280.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__1_.mem_top_track_288.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__1_.mem_top_track_288.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__1_.mem_top_track_296.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_0__1_.mem_top_track_296.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_0__1_.mem_top_track_304.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_304.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_312.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_0__1_.mem_top_track_312.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_0__1_.mem_top_track_320.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__1_.mem_top_track_320.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__1_.mem_top_track_328.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__1_.mem_top_track_328.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__1_.mem_top_track_336.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__1_.mem_top_track_336.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__1_.mem_top_track_344.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__1_.mem_top_track_344.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__1_.mem_top_track_352.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__1_.mem_top_track_352.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__1_.mem_top_track_360.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_top_track_360.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_top_track_368.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_top_track_368.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_top_track_376.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_top_track_376.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_top_track_384.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_384.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_66.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_66.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_68.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_68.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_72.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_72.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_74.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_74.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_76.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_76.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_78.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_78.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_82.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_82.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_84.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_84.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_86.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_86.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_90.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_90.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_92.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_92.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_94.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_94.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_98.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_98.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_100.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_100.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_102.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_102.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_104.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_104.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_106.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_106.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_108.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_108.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_112.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_112.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_114.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_114.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_116.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_116.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_118.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_118.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_120.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_120.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_122.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_122.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_124.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_124.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_126.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_126.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_130.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_130.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_132.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_132.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_134.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_134.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_136.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_136.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_138.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_138.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_140.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_140.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_146.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_146.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_148.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_148.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_150.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_150.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_154.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_154.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_156.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_156.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_158.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_158.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_162.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_162.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_164.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_164.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_166.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_166.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_170.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_170.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_172.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_172.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_174.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_174.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_178.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_178.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_180.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_180.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_182.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_182.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_184.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_184.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_186.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_186.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_188.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_188.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_190.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_190.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_194.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_194.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_196.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_196.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_198.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_198.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_202.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_202.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_204.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_204.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_206.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_206.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_210.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_210.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_212.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_212.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_214.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_214.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_216.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_216.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_218.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_218.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_220.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_220.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_222.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_222.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_224.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_224.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_226.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_226.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_228.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_228.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_230.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_230.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_232.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_232.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_234.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_234.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_236.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_236.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_238.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_238.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_240.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_240.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_242.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_242.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_244.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_244.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_246.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_246.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_248.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_248.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_250.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_250.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_252.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_252.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_254.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_254.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_258.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_258.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_260.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_260.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_262.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_262.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_264.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_264.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_266.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_266.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_268.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_268.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_270.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_270.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_274.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_274.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_276.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_276.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_278.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_278.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_282.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_282.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_284.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_284.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_286.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_286.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_288.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_288.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_290.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_290.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_292.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_292.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_294.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_294.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_298.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_298.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_300.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_300.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_302.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_302.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_306.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_306.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_308.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_308.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_310.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_310.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_314.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_314.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_316.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_316.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_318.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_318.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_322.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_322.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_324.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_324.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_326.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_326.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_330.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_330.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_332.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_332.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_334.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_334.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_338.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_338.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_340.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_340.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_342.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_342.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_344.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_344.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_346.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_346.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_348.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_348.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_350.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_350.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_352.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_352.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_354.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_354.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_356.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__1_.mem_right_track_356.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__1_.mem_right_track_358.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_358.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_360.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_360.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_362.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_362.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_364.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_364.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_366.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_366.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_368.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_368.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_370.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_370.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_372.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_372.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_374.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_374.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_376.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_376.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_378.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_378.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_380.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_380.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_382.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_382.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_185.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_320.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_320.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_64.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_64.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_66.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_66.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_68.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_68.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_72.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_72.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_74.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_74.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_76.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_76.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_78.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_78.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_80.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_80.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_82.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_82.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_84.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_84.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_86.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_86.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_88.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_88.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_90.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_90.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_92.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_92.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_94.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_94.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_96.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_96.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_98.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_98.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_100.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_100.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_102.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_102.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_104.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_104.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_106.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_106.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_108.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_108.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_112.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_112.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_114.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_114.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_116.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_116.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_118.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_118.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_120.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_120.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_122.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_122.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_124.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_124.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_126.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_126.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_128.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_128.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_130.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_130.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_132.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_132.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_134.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_134.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_136.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_136.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_138.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_138.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_140.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_140.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_144.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_144.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_146.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_146.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_148.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_148.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_150.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_150.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_154.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_154.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_156.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_156.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_158.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_158.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_160.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_160.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_162.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_162.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_164.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_164.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_166.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_166.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_170.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_170.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_172.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_172.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_174.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_174.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_178.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_178.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_180.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_180.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_182.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_182.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_184.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_184.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_186.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_186.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_188.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_188.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_190.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_190.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_192.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_192.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_194.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_194.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_196.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_196.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_198.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_198.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_200.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_200.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_202.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_202.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_204.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_204.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_206.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_206.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_208.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_208.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_210.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_210.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_212.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_212.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_214.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_214.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_216.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_216.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_218.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_218.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_220.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__2_.mem_right_track_220.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__2_.mem_right_track_222.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_222.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_224.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_224.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_226.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_226.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_228.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_228.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_230.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_230.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_232.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_232.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_234.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_234.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_236.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_236.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_238.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_238.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_240.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__2_.mem_right_track_240.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__2_.mem_right_track_242.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_242.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_244.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_244.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_246.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_246.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_248.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_248.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_250.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_250.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_252.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_252.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_254.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_254.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_256.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_256.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_258.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_258.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_260.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_260.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_262.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_262.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_264.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_264.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_266.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__2_.mem_right_track_266.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__2_.mem_right_track_268.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_268.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_270.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_270.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_272.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__2_.mem_right_track_272.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__2_.mem_right_track_274.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_274.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_276.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_276.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_278.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_278.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_280.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_280.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_282.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_282.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_284.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_284.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_286.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_286.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_288.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_288.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_290.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_290.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_292.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_292.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_294.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_294.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_296.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_296.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_298.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_298.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_300.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_300.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_302.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_302.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_304.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_304.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_306.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_306.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_308.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_308.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_310.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_310.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_312.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_312.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_314.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_314.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_316.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_316.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_318.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_318.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_320.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_0__2_.mem_right_track_320.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_0__2_.mem_right_track_322.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_322.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_324.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_324.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_326.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_326.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_328.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_328.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_330.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_330.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_332.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_332.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_334.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_334.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_338.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__2_.mem_right_track_338.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__2_.mem_right_track_340.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_340.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_342.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_342.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_346.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_346.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_348.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_348.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_350.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_350.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_352.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_352.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_354.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_354.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_356.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_356.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_358.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_358.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_362.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_362.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_364.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_364.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_366.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_366.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_370.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_370.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_372.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_372.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_374.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_374.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_376.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_376.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_378.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_378.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_380.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_380.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_382.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_382.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_73.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_73.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_81.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_81.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_89.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_105.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_113.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_121.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_121.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_129.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_137.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_137.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_145.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_145.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_153.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_153.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_161.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_161.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_169.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_169.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_177.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_177.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_185.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_185.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_193.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_193.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_201.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_201.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_209.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_209.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_217.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_217.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_225.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_225.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_233.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_233.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_241.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_241.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_249.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_249.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_257.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_257.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_265.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_265.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_273.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_273.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_281.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_281.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_297.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_297.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_305.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_305.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_313.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_313.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_321.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_321.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_329.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_329.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_337.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_337.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_345.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_345.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_353.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_353.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_361.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_361.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_369.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_369.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_377.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_377.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_385.mem_out[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_385.mem_outb[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_272.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_top_track_272.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_top_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_98.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_98.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_122.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_122.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_142.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_142.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_146.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_146.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_152.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_152.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_162.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_162.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_188.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_188.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_200.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_200.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_210.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_210.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_212.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_212.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_214.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_214.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_216.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_216.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_218.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_218.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_222.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_222.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_224.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_224.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_226.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_226.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_228.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_228.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_232.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_232.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_234.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_234.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_236.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_236.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_240.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_240.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_244.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_244.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_248.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_248.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_250.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_250.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_252.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_252.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_256.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_256.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_258.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_258.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_260.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_260.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_266.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_266.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_268.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_268.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_270.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_270.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_272.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_272.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_274.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_274.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_276.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_276.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_280.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_280.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_284.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_284.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_286.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_286.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_290.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_290.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_296.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_296.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_298.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_298.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_300.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_300.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_304.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_304.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_306.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_306.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_308.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_308.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_312.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_312.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_314.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_314.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_316.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_316.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_320.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_320.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_322.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_322.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_324.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_324.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_328.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_328.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_330.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_330.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_332.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_332.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_336.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_336.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_338.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_338.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_340.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_340.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_342.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_342.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_344.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_344.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_346.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_346.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_348.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_348.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_352.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_352.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_354.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_354.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_356.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_356.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_358.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_358.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_360.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_360.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_362.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_362.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_364.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_364.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_368.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_368.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_370.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_370.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_372.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_372.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_376.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_376.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_378.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_378.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_380.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_380.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_200.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_200.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_208.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_208.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_224.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_224.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_376.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_376.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_384.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_384.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_66.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_66.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_68.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_68.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_74.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_74.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_76.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_76.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_78.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_78.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_82.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_82.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_84.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_84.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_86.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_86.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_90.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_90.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_92.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_92.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_94.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_94.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_98.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_98.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_100.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_100.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_102.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_102.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_106.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_106.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_108.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_108.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_114.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_114.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_116.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_116.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_118.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_118.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_122.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_122.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_124.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_124.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_126.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_126.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_130.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_130.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_132.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_132.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_134.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_134.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_138.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_138.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_140.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_140.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_146.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_146.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_148.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_148.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_150.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_150.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_154.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_154.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_156.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_156.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_158.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_158.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_162.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_162.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_164.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_164.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_166.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_166.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_168.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_168.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_170.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_170.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_172.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_172.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_174.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_174.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_178.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_178.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_180.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_180.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_182.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_182.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_186.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_186.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_188.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_188.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_190.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_190.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_192.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_192.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_194.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_194.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_196.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_196.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_198.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_198.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_202.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_202.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_204.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_204.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_206.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_206.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_210.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_210.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_212.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_212.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_214.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_214.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_218.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_218.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_220.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_220.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_222.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_222.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_226.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_226.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_228.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_228.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_230.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_230.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_234.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_234.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_236.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_236.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_238.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_238.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_242.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_242.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_244.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_244.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_246.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_246.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_250.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_250.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_252.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_252.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_254.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_254.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_258.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_258.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_260.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_260.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_262.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_262.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_266.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_266.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_268.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_268.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_270.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_270.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_274.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_274.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_276.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_276.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_278.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_278.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_282.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_282.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_284.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_284.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_286.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_286.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_290.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_290.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_292.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_292.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_294.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_294.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_298.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_298.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_300.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_300.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_302.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_302.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_306.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_306.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_308.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_308.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_310.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_310.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_314.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_314.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_316.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_316.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_318.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_318.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_322.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_322.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_324.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_324.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_326.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_326.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_330.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_330.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_332.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_332.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_334.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_334.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_338.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_338.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_340.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_340.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_342.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_342.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_346.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_346.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_348.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_348.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_350.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_350.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_354.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_354.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_356.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_356.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_358.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_358.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_362.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_362.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_364.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_364.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_366.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_366.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_370.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_370.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_372.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_372.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_374.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_374.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_376.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_376.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_378.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_378.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_380.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_380.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_382.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_382.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_66.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_66.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_68.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_68.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_74.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_74.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_76.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_76.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_78.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_78.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_82.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_82.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_84.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_84.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_86.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_86.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_90.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_90.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_92.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_92.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_94.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_94.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_98.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_98.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_100.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_100.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_102.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_102.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_106.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_106.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_108.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_108.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_114.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_114.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_116.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_116.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_118.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_118.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_122.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_122.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_124.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_124.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_126.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_126.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_130.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_130.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_132.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_132.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_134.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_134.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_138.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_138.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_140.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_140.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_146.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_146.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_148.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_148.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_150.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_150.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_154.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_154.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_156.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_156.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_158.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_158.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_162.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_162.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_164.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_164.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_166.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_166.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_170.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_170.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_172.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_172.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_174.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_174.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_178.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_178.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_180.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_180.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_182.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_182.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_186.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_186.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_188.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_188.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_190.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_190.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_194.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_194.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_196.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_196.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_198.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_198.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_202.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_202.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_204.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_204.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_206.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_206.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_210.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_210.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_212.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_212.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_214.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_214.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_218.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_218.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_220.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_220.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_222.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_222.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_226.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_226.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_228.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_228.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_230.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_230.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_234.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_234.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_236.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_236.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_238.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_238.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_242.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_242.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_244.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_244.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_246.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_246.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_250.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_250.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_252.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_252.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_254.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_254.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_258.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_258.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_260.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_260.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_262.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_262.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_266.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_266.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_268.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_268.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_270.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_270.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_274.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_274.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_276.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_276.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_278.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_278.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_282.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_282.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_284.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_284.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_286.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_286.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_290.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_290.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_292.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_292.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_294.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_294.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_298.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_298.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_300.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_300.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_302.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_302.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_306.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_306.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_308.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_308.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_310.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_310.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_314.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_314.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_316.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_316.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_318.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_318.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_322.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_322.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_324.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_324.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_326.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_326.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_330.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_330.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_332.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_332.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_334.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_334.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_336.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_336.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_338.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_338.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_340.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_340.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_342.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_342.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_346.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_346.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_348.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_348.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_350.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_350.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_354.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_354.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_356.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_356.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_358.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_358.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_360.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_360.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_362.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_362.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_364.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_364.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_366.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_366.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_370.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_370.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_372.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_372.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_374.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_374.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_376.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_376.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_378.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_378.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_380.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_380.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_382.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_382.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_113.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_113.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_193.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_193.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_201.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_201.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_321.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_321.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_337.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_337.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_361.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_361.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_369.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_369.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_377.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_377.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_210.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_210.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_212.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_212.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_216.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_216.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_218.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_218.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_222.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_222.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_224.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_224.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_226.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_226.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_228.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_228.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_234.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_234.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_236.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_236.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_240.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_240.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_244.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_244.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_248.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_248.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_252.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_252.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_256.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_256.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_258.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_258.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_260.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_260.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_266.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_266.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_270.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_270.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_272.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_272.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_274.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_274.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_276.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_276.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_280.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_280.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_284.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_284.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_288.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_288.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_290.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_290.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_296.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_296.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_298.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_298.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_300.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_300.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_306.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_306.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_308.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_308.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_312.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_312.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_314.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_314.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_316.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_316.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_320.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_320.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_324.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_324.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_328.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_328.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_330.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_330.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_332.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_332.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_336.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_336.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_338.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_338.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_342.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_342.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_344.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_344.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_346.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_346.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_348.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_348.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_352.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_352.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_354.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_354.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_356.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_356.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_360.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_360.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_362.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_362.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_364.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_364.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_368.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_368.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_370.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_370.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_372.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_372.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_376.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_376.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_378.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_378.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_380.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_380.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_384.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_384.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_215.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_215.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_233.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_233.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_251.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_251.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_269.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_269.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_287.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_287.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_305.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_305.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_323.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_323.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_341.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_341.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_359.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_359.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_100.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_100.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_106.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_106.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_130.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_130.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_148.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_148.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_152.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_152.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_154.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_154.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_190.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_190.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_202.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_202.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_208.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_208.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_210.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_210.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_212.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_212.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_214.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_214.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_216.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_216.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_218.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_218.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_222.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_222.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_224.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_224.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_226.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_226.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_228.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_228.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_232.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_232.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_234.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_234.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_236.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_236.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_240.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_240.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_244.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_244.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_248.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_248.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_250.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_250.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_252.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_252.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_256.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_256.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_258.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_258.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_260.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_260.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_266.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_266.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_268.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_268.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_270.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_270.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_272.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_272.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_274.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_274.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_276.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_276.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_280.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_280.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_284.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_284.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_290.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_290.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_296.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_296.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_298.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_298.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_300.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_300.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_304.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_304.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_306.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_306.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_308.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_308.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_312.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_312.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_314.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_314.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_316.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_316.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_320.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_320.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_322.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_322.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_324.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_324.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_328.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_328.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_330.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_330.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_332.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_332.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_336.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_336.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_338.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_338.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_340.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_340.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_342.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_342.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_344.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_344.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_346.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_346.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_348.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_348.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_352.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_352.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_354.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_354.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_356.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_356.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_358.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_358.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_360.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_360.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_362.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_362.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_364.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_364.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_368.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_368.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_370.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_370.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_372.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_372.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_376.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_376.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_378.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_378.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_380.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_380.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_136.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_136.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_144.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_144.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_152.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_152.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_160.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_right_track_160.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_192.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_192.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_208.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_208.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_232.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_232.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_240.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_240.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_256.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_right_track_256.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_right_track_264.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_264.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_272.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_272.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_296.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_296.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_304.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_304.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_312.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_right_track_312.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_right_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_328.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_328.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_344.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_344.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_352.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_352.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_360.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_360.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_376.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_376.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__1_.mem_top_track_72.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_72.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_80.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__1_.mem_top_track_80.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__1_.mem_top_track_88.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_top_track_88.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_top_track_96.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_96.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_104.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_1__1_.mem_top_track_104.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_1__1_.mem_top_track_112.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__1_.mem_top_track_112.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__1_.mem_top_track_120.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_120.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_128.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_top_track_128.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_top_track_136.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__1_.mem_top_track_136.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__1_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_152.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_top_track_152.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_top_track_160.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_top_track_160.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_top_track_168.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_top_track_168.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_top_track_176.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_top_track_176.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_top_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_192.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__1_.mem_top_track_192.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__1_.mem_top_track_200.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_1__1_.mem_top_track_200.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_1__1_.mem_top_track_208.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_208.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_216.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__1_.mem_top_track_216.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__1_.mem_top_track_224.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_1__1_.mem_top_track_224.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_1__1_.mem_top_track_232.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_232.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_248.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_top_track_248.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_top_track_256.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_top_track_256.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_top_track_264.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__1_.mem_top_track_264.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__1_.mem_top_track_272.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_top_track_272.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_top_track_280.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_top_track_280.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_top_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_296.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_296.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_304.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__1_.mem_top_track_304.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__1_.mem_top_track_312.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__1_.mem_top_track_312.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__1_.mem_top_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_336.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__1_.mem_top_track_336.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__1_.mem_top_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_352.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_352.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_360.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_top_track_360.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_top_track_368.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__1_.mem_top_track_368.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__1_.mem_top_track_376.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_376.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_384.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__1_.mem_top_track_384.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_80.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_88.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_88.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_96.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_96.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_104.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_112.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_112.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_128.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_136.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_136.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_144.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_144.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_152.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_160.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_160.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_176.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_184.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_184.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_192.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__1_.mem_right_track_192.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__1_.mem_right_track_200.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_216.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__1_.mem_right_track_216.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__1_.mem_right_track_224.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_224.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_232.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_232.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_240.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__1_.mem_right_track_240.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__1_.mem_right_track_248.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_248.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_256.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_256.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_264.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__1_.mem_right_track_264.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__1_.mem_right_track_272.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_272.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_280.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_280.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_288.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__1_.mem_right_track_288.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__1_.mem_right_track_296.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_296.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_304.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_304.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_320.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_320.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_328.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_328.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_336.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__1_.mem_right_track_336.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__1_.mem_right_track_344.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_344.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_360.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__1_.mem_right_track_360.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__1_.mem_right_track_368.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_368.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_384.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__1_.mem_right_track_384.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_105.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_105.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_145.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_145.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_185.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_185.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_273.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_273.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_289.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_289.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_305.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_305.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_329.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_329.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_345.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_345.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_353.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_353.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_361.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_361.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_369.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_369.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_193.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_left_track_193.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_left_track_201.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_201.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_217.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_217.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_321.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_321.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_337.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_337.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_361.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_361.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_369.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_369.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_377.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_377.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_112.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_top_track_112.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_272.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_top_track_272.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_312.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_top_track_312.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_376.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__2_.mem_top_track_376.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__2_.mem_top_track_384.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__2_.mem_top_track_384.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_80.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_right_track_80.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_right_track_88.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__2_.mem_right_track_88.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__2_.mem_right_track_96.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_96.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_104.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__2_.mem_right_track_104.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__2_.mem_right_track_112.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_112.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_120.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__2_.mem_right_track_120.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__2_.mem_right_track_128.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__2_.mem_right_track_128.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__2_.mem_right_track_136.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_right_track_136.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_152.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_right_track_152.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_184.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_184.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_192.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_192.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_208.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__2_.mem_right_track_208.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__2_.mem_right_track_216.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__2_.mem_right_track_216.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__2_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_232.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_right_track_232.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_248.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_248.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_256.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_256.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_280.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_right_track_280.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_296.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_296.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_304.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__2_.mem_right_track_304.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__2_.mem_right_track_312.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_312.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_320.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_320.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_328.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_328.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_344.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__2_.mem_right_track_344.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__2_.mem_right_track_352.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__2_.mem_right_track_352.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__2_.mem_right_track_360.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_360.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_368.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_368.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_384.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_1__2_.mem_right_track_384.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_73.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_73.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_81.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_81.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_89.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_97.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_97.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_105.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_113.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_121.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_121.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_129.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_137.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_137.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_145.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_145.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_153.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_153.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_161.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_161.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_169.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_169.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_177.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_177.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_185.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_185.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_193.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_193.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_201.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_201.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_209.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_209.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_217.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_217.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_225.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_225.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_233.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_233.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_241.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_241.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_249.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_249.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_257.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_257.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_265.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_265.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_273.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_273.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_281.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_281.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_289.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_289.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_297.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_297.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_305.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_305.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_313.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_313.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_321.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_321.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_329.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_329.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_337.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_337.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_345.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_345.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_353.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_353.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_361.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_361.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_369.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_369.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_377.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_377.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_385.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_385.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_193.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_193.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_201.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_201.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_321.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_321.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_337.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_337.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_361.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_361.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_369.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_369.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_377.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_377.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_80.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_80.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_88.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_right_track_88.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_right_track_96.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_96.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_104.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_104.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_136.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_right_track_136.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_152.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_152.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_216.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_216.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_224.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_224.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_248.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_248.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_256.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_right_track_256.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_right_track_264.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_264.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_272.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_272.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_280.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_right_track_280.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_296.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_296.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_344.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_344.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_360.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_360.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_368.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__3_.mem_right_track_368.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__3_.mem_right_track_376.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_1__3_.mem_right_track_376.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_1__3_.mem_right_track_384.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_1__3_.mem_right_track_384.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_81.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_81.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_129.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_129.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_169.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_169.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_289.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_289.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_361.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_361.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_385.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_385.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_200.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_200.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_208.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_208.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_224.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_224.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_360.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_360.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_368.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_368.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_376.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_376.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_384.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_384.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_72.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__4_.mem_right_track_72.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_104.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__4_.mem_right_track_104.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_120.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__4_.mem_right_track_120.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_136.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__4_.mem_right_track_136.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_168.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__4_.mem_right_track_168.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_216.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__4_.mem_right_track_216.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__4_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_320.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__4_.mem_right_track_320.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__4_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_273.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_273.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_329.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_329.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_361.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_361.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_193.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_193.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_201.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_201.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_321.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_321.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_337.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_337.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_361.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_361.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_369.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_369.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_377.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_377.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_72.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__5_.mem_right_track_72.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_176.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__5_.mem_right_track_176.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_200.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__5_.mem_right_track_200.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__5_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_264.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__5_.mem_right_track_264.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__5_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_360.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__5_.mem_right_track_360.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__5_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_193.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_193.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_201.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_201.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_289.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_289.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_297.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_297.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_321.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_321.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_337.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_337.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_361.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_361.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_369.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_369.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_377.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_377.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_193.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_193.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_201.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_201.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_321.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_321.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_337.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_337.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_361.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__5_.mem_left_track_361.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__5_.mem_left_track_369.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_369.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_377.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_377.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_215.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_215.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_217.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_217.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_233.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_233.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_235.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_235.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_251.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_251.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_253.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_253.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_269.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_269.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_271.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_271.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_287.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_287.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_289.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_289.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_305.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_305.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_307.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_307.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_323.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_323.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_325.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_325.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_341.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_341.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_343.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_343.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_359.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_359.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_379.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_379.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_104.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_104.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_152.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_152.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_194.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_194.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_210.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_210.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_212.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_212.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_214.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_214.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_216.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_216.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_218.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_218.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_222.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_222.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_224.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_224.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_226.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_226.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_228.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_228.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_232.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_232.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_234.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_234.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_236.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_236.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_240.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_240.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_244.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_244.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_248.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_248.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_250.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_250.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_252.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_252.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_256.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_256.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_258.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_258.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_260.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_260.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_266.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_266.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_268.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_268.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_270.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_270.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_272.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_272.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_274.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_274.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_276.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_276.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_280.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_280.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_284.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_284.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_290.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_290.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_296.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_296.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_298.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_298.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_300.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_300.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_304.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_304.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_306.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_306.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_308.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_308.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_312.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_312.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_314.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_314.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_316.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_316.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_320.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_320.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_322.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_322.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_324.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_324.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_328.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_328.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_330.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_330.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_332.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_332.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_336.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_336.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_338.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_338.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_340.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_340.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_342.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_342.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_344.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_344.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_346.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_346.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_348.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_348.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_352.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_352.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_354.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_354.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_356.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_356.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_358.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_358.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_360.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_360.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_362.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_362.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_364.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_364.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_368.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_368.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_370.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_370.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_372.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_372.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_376.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_376.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_378.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_378.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_380.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_380.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_72.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_72.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_80.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_88.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_right_track_88.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_right_track_96.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_96.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_104.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_104.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_112.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_120.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_120.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_128.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_128.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_136.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_152.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_right_track_152.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_right_track_160.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_160.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_200.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_200.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_216.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_216.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_224.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_224.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_232.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_232.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_240.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_240.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_248.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_248.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_256.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_256.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_264.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_264.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_272.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_272.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_280.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_right_track_280.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_right_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_304.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_304.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_312.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_312.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_320.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_320.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_336.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_336.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_352.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_352.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_360.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_360.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_368.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_368.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_72.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_72.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_80.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_80.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_104.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_104.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_192.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_192.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_200.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_200.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_232.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_232.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_240.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_240.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_248.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_248.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_256.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_256.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_272.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_top_track_272.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_288.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_288.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_296.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_296.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_304.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_304.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_320.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_320.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_344.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_344.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_368.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_368.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_384.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_top_track_384.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_88.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_88.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_96.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_96.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_104.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_128.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_136.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_right_track_136.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_right_track_144.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_144.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_168.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_168.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_184.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_right_track_184.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_right_track_192.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_right_track_192.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_216.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_right_track_216.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_232.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_232.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_256.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_right_track_256.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_right_track_264.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_264.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_296.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_right_track_296.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_right_track_304.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_right_track_304.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_320.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_right_track_320.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_336.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_right_track_336.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_right_track_344.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_right_track_344.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_right_track_352.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_352.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_360.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_360.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_177.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_177.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_225.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_225.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_249.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_249.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_257.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_257.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_273.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_273.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_208.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_top_track_208.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_top_track_216.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_216.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_224.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_top_track_224.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_248.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_top_track_248.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_296.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_top_track_296.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_72.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_right_track_72.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_right_track_80.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_80.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_88.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_88.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_96.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_96.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_104.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_120.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_120.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_144.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_144.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_152.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_right_track_152.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_right_track_160.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_160.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_168.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_right_track_168.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_184.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__2_.mem_right_track_184.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__2_.mem_right_track_192.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_192.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_200.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_200.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_224.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_right_track_224.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_right_track_232.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_232.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_240.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_240.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_248.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_248.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_256.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_256.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_264.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_264.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_280.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__2_.mem_right_track_280.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__2_.mem_right_track_288.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_288.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_304.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_right_track_304.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_320.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_320.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_328.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__2_.mem_right_track_328.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__2_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_344.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_344.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_352.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_right_track_352.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_368.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_right_track_368.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_right_track_376.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_right_track_376.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_right_track_384.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_right_track_384.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_73.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_73.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_81.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_81.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_89.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_89.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_121.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_121.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_145.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_145.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_153.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_153.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_161.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_161.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_185.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_185.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_193.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_193.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_201.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_201.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_209.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_209.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_217.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_217.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_225.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_225.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_233.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_233.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_241.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_241.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_249.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_249.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_257.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_257.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_281.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_281.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_289.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_289.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_297.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_297.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_305.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_305.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_313.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_313.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_329.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_329.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_337.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_337.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_345.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_345.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_361.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_361.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_377.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_377.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_385.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_left_track_385.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_160.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__3_.mem_top_track_160.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_120.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_right_track_120.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_right_track_128.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_right_track_128.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_144.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_144.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_152.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_right_track_152.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_176.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_right_track_176.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_right_track_184.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_184.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_352.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_352.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_105.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_105.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_233.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_233.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_289.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_289.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_305.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_305.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_313.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_313.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_321.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_321.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_345.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_345.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_353.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_353.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_369.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_369.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_377.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_377.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_265.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_left_track_265.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_256.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_right_track_256.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_right_track_264.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__4_.mem_right_track_264.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__4_.mem_right_track_272.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__4_.mem_right_track_272.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__4_.mem_right_track_280.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_right_track_280.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_right_track_288.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__4_.mem_right_track_288.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__4_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_312.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__4_.mem_right_track_312.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__4_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_376.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__4_.mem_right_track_376.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__4_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_281.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_281.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_80.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_right_track_80.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_280.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_right_track_280.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_336.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_right_track_336.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_89.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_89.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_129.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_129.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_209.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_209.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_289.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_289.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_305.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_305.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_329.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_329.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_215.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_215.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_217.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_217.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_233.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_233.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_235.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_235.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_251.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_251.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_253.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_253.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_269.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_269.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_271.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_271.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_287.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_287.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_289.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_289.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_305.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_305.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_307.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_307.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_323.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_323.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_325.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_325.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_341.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_341.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_343.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_343.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_359.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_359.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_379.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_379.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_114.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_114.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_120.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_120.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_126.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_126.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_138.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_138.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_146.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_146.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_152.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_152.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_156.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_156.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_160.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_160.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_162.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_162.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_178.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_178.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_180.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_180.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_184.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_184.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_186.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_186.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_198.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_198.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_200.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_200.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_202.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_202.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_204.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_204.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_210.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_210.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_212.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_212.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_214.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_214.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_216.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_216.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_218.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_218.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_222.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_222.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_224.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_224.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_226.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_226.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_228.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_228.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_232.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_232.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_234.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_234.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_236.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_236.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_240.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_240.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_244.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_244.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_248.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_248.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_250.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_250.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_252.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_252.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_256.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_256.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_258.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_258.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_260.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_260.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_266.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_266.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_268.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_268.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_270.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_270.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_272.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_272.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_274.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_274.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_276.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_276.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_280.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_280.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_284.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_284.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_290.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_290.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_296.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_296.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_298.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_298.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_300.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_300.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_304.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_304.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_306.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_306.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_308.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_308.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_312.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_312.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_314.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_314.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_316.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_316.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_320.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_320.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_322.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_322.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_324.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_324.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_328.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_328.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_330.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_330.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_332.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_332.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_336.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_336.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_338.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_338.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_340.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_340.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_342.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_342.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_344.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_344.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_346.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_346.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_348.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_348.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_352.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_352.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_354.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_354.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_356.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_356.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_358.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_358.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_360.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_360.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_362.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_362.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_364.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_364.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_368.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_368.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_370.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_370.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_372.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_372.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_376.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_376.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_378.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_378.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_380.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_380.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_72.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_72.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_88.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_88.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_120.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_120.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_128.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_right_track_128.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_right_track_136.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_136.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_152.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_152.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_168.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_168.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_184.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_184.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_208.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_208.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_224.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_right_track_224.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_right_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_248.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_248.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_272.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_272.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_312.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_312.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_72.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_72.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_80.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_top_track_80.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_top_track_88.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_88.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_104.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_top_track_104.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_top_track_112.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_112.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_120.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_120.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_128.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_top_track_128.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_top_track_136.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_136.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_144.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_144.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_152.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_152.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_160.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_160.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_168.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_168.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_176.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_176.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_184.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_184.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_192.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_192.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_200.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_200.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_208.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_208.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_216.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_216.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_224.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_224.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_232.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_232.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_240.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_240.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_248.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_248.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_256.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_256.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_264.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_264.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_272.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_272.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_280.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_280.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_288.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_288.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_296.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_top_track_296.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_top_track_304.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_304.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_312.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_312.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_320.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_320.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_328.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_328.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_336.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_336.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_344.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_344.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_352.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_352.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_360.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_360.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_top_track_368.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_top_track_368.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_top_track_376.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_376.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_384.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_384.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_72.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_right_track_72.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_right_track_80.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_80.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_96.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__1_.mem_right_track_96.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__1_.mem_right_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_120.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_right_track_120.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_right_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_144.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_right_track_144.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_right_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_160.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_160.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_168.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_right_track_168.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_right_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_200.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_200.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_208.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_208.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_216.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_right_track_216.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_right_track_224.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_224.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_232.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_232.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_256.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_right_track_256.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_right_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_272.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_272.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_312.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_312.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_320.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__1_.mem_right_track_320.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__1_.mem_right_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_360.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_360.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_368.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_368.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_376.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_376.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_384.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_384.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_88.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_88.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_120.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__2_.mem_right_track_120.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__2_.mem_right_track_128.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_right_track_128.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_right_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_152.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__2_.mem_right_track_152.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__2_.mem_right_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_168.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_168.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_192.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__2_.mem_right_track_192.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__2_.mem_right_track_200.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__2_.mem_right_track_200.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__2_.mem_right_track_208.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__2_.mem_right_track_208.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__2_.mem_right_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_224.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__2_.mem_right_track_224.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__2_.mem_right_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_240.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__2_.mem_right_track_240.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__2_.mem_right_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_264.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__2_.mem_right_track_264.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__2_.mem_right_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_328.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_328.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_344.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_right_track_344.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_right_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_360.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_360.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_368.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__2_.mem_right_track_368.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__2_.mem_right_track_376.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_376.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_384.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_384.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_73.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_73.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_89.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_105.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_113.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_129.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_137.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_137.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_153.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_153.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_169.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_169.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_177.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_177.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_185.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_185.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_193.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_193.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_201.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_201.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_225.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_225.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_233.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_233.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_241.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_241.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_249.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_249.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_257.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_257.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_273.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_273.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_297.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_297.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_313.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_313.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_321.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_321.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_329.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_329.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_337.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_337.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_345.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_345.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_353.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_353.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_361.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_361.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_369.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_369.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_377.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_377.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_313.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_313.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_73.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_73.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_129.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_129.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_137.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_137.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_153.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_153.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_161.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_161.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_193.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_193.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_209.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_209.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_217.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_217.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_257.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_257.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_265.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_265.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_289.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_289.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_329.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_329.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_353.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_353.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_377.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_377.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_113.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__3_.mem_left_track_113.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_200.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_200.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_208.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_208.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_224.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_224.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_360.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_360.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_368.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_368.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_376.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_376.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_384.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_384.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_200.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_200.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_208.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_208.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_224.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_224.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_360.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_360.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_368.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_368.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_376.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_376.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_384.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_384.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_73.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_73.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_105.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_105.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_121.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_121.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_145.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_145.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_177.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_177.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_193.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_193.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_201.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_201.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_273.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_273.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_297.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_297.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_321.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_321.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_337.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_337.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_361.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_361.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_369.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_369.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_152.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_152.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_160.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_160.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_168.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_168.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_176.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_176.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_184.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_184.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_192.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_192.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_200.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_200.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_208.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_208.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_216.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_216.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_224.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_224.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_232.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_232.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_240.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_240.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_248.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_248.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_256.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_256.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_264.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_264.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_272.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_272.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_280.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_280.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_288.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_288.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_296.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_296.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_304.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_304.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_312.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_312.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_320.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_320.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_328.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_328.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_336.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_336.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_344.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_344.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_352.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_352.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_360.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_360.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_368.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_368.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_384.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_384.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_200.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_200.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_208.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_208.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_224.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_224.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_360.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_360.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_368.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_368.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_376.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_376.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_384.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_384.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_193.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_193.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_201.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_201.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_209.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_209.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_217.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_217.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_305.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_305.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_321.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_321.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_337.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_337.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_353.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_353.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_361.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_361.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_369.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_369.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_377.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_377.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_215.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_215.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_217.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_217.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_233.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_233.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_235.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_235.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_251.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_251.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_253.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_253.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_269.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_269.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_271.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_271.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_287.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_287.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_289.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_289.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_305.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_305.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_307.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_307.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_323.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_323.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_325.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_325.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_341.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_341.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_343.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_343.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_359.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_359.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_379.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_379.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_74.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_74.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_80.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_80.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_86.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_86.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_104.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_104.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_106.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_106.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_112.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_112.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_114.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_114.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_120.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_120.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_128.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_128.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_138.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_138.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_146.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_146.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_148.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_148.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_150.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_150.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_152.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_152.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_154.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_154.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_156.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_156.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_158.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_158.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_160.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_160.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_164.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_164.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_166.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_166.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_168.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_168.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_170.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_170.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_172.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_172.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_174.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_174.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_176.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_176.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_178.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_178.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_180.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_180.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_182.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_182.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_184.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_184.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_186.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_186.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_188.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_188.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_190.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_190.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_192.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_192.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_194.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_194.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_196.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_196.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_200.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_200.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_202.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_202.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_204.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_204.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_206.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_206.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_208.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_208.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_210.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_210.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_212.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_212.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_214.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_214.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_218.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_218.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_220.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_220.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_222.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_222.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_224.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_224.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_226.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_226.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_228.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_228.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_230.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_230.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_232.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_232.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_236.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_236.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_238.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_238.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_240.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_240.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_242.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_242.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_244.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_244.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_246.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_246.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_248.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_248.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_250.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_250.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_254.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_254.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_256.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_256.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_258.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_258.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_260.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_260.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_262.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_262.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_264.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_264.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_266.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_266.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_268.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_268.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_272.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_272.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_274.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_274.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_276.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_276.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_278.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_278.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_280.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_280.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_282.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_282.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_284.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_284.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_286.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_286.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_290.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_290.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_292.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_292.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_294.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_294.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_296.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_296.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_298.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_298.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_300.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_300.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_302.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_302.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_304.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_304.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_308.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_308.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_310.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_310.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_312.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_312.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_314.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_314.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_316.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_316.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_318.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_318.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_320.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_320.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_322.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_322.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_326.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_326.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_328.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_328.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_330.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_330.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_332.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_332.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_334.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_334.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_336.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_336.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_338.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_338.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_340.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_340.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_344.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_344.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_346.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_346.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_348.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_348.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_350.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_350.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_352.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_352.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_354.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_354.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_356.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_356.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_358.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_358.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_360.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_360.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_362.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_362.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_364.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_364.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_366.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_366.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_368.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_368.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_370.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_370.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_372.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_372.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_374.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_374.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_376.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_376.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_380.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_380.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_382.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_382.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_384.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_384.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_215.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_215.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_217.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_217.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_233.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_233.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_235.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_235.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_251.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_251.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_253.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_253.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_269.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_269.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_271.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_271.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_287.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_287.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_289.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_289.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_305.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_305.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_307.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_307.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_323.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_323.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_325.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_325.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_341.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_341.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_343.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_343.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_359.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_359.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_379.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_379.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_72.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__1_.mem_top_track_72.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__1_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_88.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__1_.mem_top_track_88.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__1_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_112.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__1_.mem_top_track_112.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__1_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_144.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__1_.mem_top_track_144.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__1_.mem_top_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_200.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_200.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_208.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_208.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_224.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_224.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_240.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__1_.mem_top_track_240.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__1_.mem_top_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_280.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__1_.mem_top_track_280.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__1_.mem_top_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_352.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__1_.mem_top_track_352.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__1_.mem_top_track_360.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__1_.mem_top_track_360.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__1_.mem_top_track_368.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_368.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_376.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_376.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_384.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_384.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_21.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_23.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_left_track_23.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_27.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_27.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_35.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_35.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_53.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_53.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_67.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_67.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_69.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_69.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_83.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_83.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_85.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_85.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_99.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_99.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_101.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_101.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_103.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_103.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_107.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_107.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_115.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_115.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_127.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_127.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_133.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_133.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_139.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_139.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_147.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_147.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_149.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_149.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_151.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_151.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_155.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_155.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_157.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_157.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_159.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_159.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_163.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_163.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_165.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_165.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_167.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_167.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_171.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_171.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_173.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_173.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_175.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_175.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_179.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_179.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_181.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_181.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_183.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_183.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_187.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_187.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_189.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_189.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_191.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_191.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_195.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_195.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_197.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_197.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_199.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_199.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_203.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_203.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_205.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_205.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_207.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_207.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_211.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_211.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_213.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_213.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_215.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_215.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_219.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_219.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_221.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_221.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_223.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_223.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_227.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_227.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_229.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_229.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_231.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_231.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_235.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_235.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_237.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_237.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_239.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_239.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_243.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_243.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_245.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_245.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_247.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_247.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_251.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_251.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_253.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_253.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_255.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_255.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_259.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_259.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_261.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_261.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_263.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_263.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_267.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_267.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_269.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_269.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_271.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_271.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_275.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_275.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_277.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_277.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_279.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_279.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_283.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_283.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_285.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_285.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_287.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_287.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_291.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_291.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_293.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_293.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_295.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_295.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_299.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_299.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_301.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_301.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_303.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_303.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_307.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_307.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_309.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_309.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_311.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_311.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_315.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_315.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_317.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_317.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_319.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_319.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_323.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_323.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_325.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_325.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_327.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_327.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_331.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_331.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_333.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_333.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_335.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_335.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_339.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_339.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_341.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_341.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_343.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_343.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_347.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_347.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_349.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_349.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_351.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_351.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_355.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_355.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_357.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_357.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_359.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_359.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_363.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_363.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_365.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_365.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_367.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_367.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_369.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_left_track_369.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_left_track_371.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_371.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_373.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_373.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_375.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_375.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_377.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_377.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_379.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_379.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_381.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_381.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_383.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_383.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_81.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_81.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_89.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_97.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_97.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_105.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_113.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_121.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_121.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_129.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_145.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_145.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_177.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_177.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_185.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_185.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_193.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_193.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_201.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_201.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_209.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_209.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_225.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_225.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_233.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_233.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_241.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_241.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_257.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_257.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_273.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_273.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_281.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_281.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_289.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_289.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_305.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_305.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_321.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_321.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_337.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_337.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_369.mem_out[0:3] = 4'b1100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_369.mem_outb[0:3] = 4'b0011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_377.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_377.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_385.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_385.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_21.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_27.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_27.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_35.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_35.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_53.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_53.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_67.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_67.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_69.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_69.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_83.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_83.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_85.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_85.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_99.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__2_.mem_left_track_99.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__2_.mem_left_track_101.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_101.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_103.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_103.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_107.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_107.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_139.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_139.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_147.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_147.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_149.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_149.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_151.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_151.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_155.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_155.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_157.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_157.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_159.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_159.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_163.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_163.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_165.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_165.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_167.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_167.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_171.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_171.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_173.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_173.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_175.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_175.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_179.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_179.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_181.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_181.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_183.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_183.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_187.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_187.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_189.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_189.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_191.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_191.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_195.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_195.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_197.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_197.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_199.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_199.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_203.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_203.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_205.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_205.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_207.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_207.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_211.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_211.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_213.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_213.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_215.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_215.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_219.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_219.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_221.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_221.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_223.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_223.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_227.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_227.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_229.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_229.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_231.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_231.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_235.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_235.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_237.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_237.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_239.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_239.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_243.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_243.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_245.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_245.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_247.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_247.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_251.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_251.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_253.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_253.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_255.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_255.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_259.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_259.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_261.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_261.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_263.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_263.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_267.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_267.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_269.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_269.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_271.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_271.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_275.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_275.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_277.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_277.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_279.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_279.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_283.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_283.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_285.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_285.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_287.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_287.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_291.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_291.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_293.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_293.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_295.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_295.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_299.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_299.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_301.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_301.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_303.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_303.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_307.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_307.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_309.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_309.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_311.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_311.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_315.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_315.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_317.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_317.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_319.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_319.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_323.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_323.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_325.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_325.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_327.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_327.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_331.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_331.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_333.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_333.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_335.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_335.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_339.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_339.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_341.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_341.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_343.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_343.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_347.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_347.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_349.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_349.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_351.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_351.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_355.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_355.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_357.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_357.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_359.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_359.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_363.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_363.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_365.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_365.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_367.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_367.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_371.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_371.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_373.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_373.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_375.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_375.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_377.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_377.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_379.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_379.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_381.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_381.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_383.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_383.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_121.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_121.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_137.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_137.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_161.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_161.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_185.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_185.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_209.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_209.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_233.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_233.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_249.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_249.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_281.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_281.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_289.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_289.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_297.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_297.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_313.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_313.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_337.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_337.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_345.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_345.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_361.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_361.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_161.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_161.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_163.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_163.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_179.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_179.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_215.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_215.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_217.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_217.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_233.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_233.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_235.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_235.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_251.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_251.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_253.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_253.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_269.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_269.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_271.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_271.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_287.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_287.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_289.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_289.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_305.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_305.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_307.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_307.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_323.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_323.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_325.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_325.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_341.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_341.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_343.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_343.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_359.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_359.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_379.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_379.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_152.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_152.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_160.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_160.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_168.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_168.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_176.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_176.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_184.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_184.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_192.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_192.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_200.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_200.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_208.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_208.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_216.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_216.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_224.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_224.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_232.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_232.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_240.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_240.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_248.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_248.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_256.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_256.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_264.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_264.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_272.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_272.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_280.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_280.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_288.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_288.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_296.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_296.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_304.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_304.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_312.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_312.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_320.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_320.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_328.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_328.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_336.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_336.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_344.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_344.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_352.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_352.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_360.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_360.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_368.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_368.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_376.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_376.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_384.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_384.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_89.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_89.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_153.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_153.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_161.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_161.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_169.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_169.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_177.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_177.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_185.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_185.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_193.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_193.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_201.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_201.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_209.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_209.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_217.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_217.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_225.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_225.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_233.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_233.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_241.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_241.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_249.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_249.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_257.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_257.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_265.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_265.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_273.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_273.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_281.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_281.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_289.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_289.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_297.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_297.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_305.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_305.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_313.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_313.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_321.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_321.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_329.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_329.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_337.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_337.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_345.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_345.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_353.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_353.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_361.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_361.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_369.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_369.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_377.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_377.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_385.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_385.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_21.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_27.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_27.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_35.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_35.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_53.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_53.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_67.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_67.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_69.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_69.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_83.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_83.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_85.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_85.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_99.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_99.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_101.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_101.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_103.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_103.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_107.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_107.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_139.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_139.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_147.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_147.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_149.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_149.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_151.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_151.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_155.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_155.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_157.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_157.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_159.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_159.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_163.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_163.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_165.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_165.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_167.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_167.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_171.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_171.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_173.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_173.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_175.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_175.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_179.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_179.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_181.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_181.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_183.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_183.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_187.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_187.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_189.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_189.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_191.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_191.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_195.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_195.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_197.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_197.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_199.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_199.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_203.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_203.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_205.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_205.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_207.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_207.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_211.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_211.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_213.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_213.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_215.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_215.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_219.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_219.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_221.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_221.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_223.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_223.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_227.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_227.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_229.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_229.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_231.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_231.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_235.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_235.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_237.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_237.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_239.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_239.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_243.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_243.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_245.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_245.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_247.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_247.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_251.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_251.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_253.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_253.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_255.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_255.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_259.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_259.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_261.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_261.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_263.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_263.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_267.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_267.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_269.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_269.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_271.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_271.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_275.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_275.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_277.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_277.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_279.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_279.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_283.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_283.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_285.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_285.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_287.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_287.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_291.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_291.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_293.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_293.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_295.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_295.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_299.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_299.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_301.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_301.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_303.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_303.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_307.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_307.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_309.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_309.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_311.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_311.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_315.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_315.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_317.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_317.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_319.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_319.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_323.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_323.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_325.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_325.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_327.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_327.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_331.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_331.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_333.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_333.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_335.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_335.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_339.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_339.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_341.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_341.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_343.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_343.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_347.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_347.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_349.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_349.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_351.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_351.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_355.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_355.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_357.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_357.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_359.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_359.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_363.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_363.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_365.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_365.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_367.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_367.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_371.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_371.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_373.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_373.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_375.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_375.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_377.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_377.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_379.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_379.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_381.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_381.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_383.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_383.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_152.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_152.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_160.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_160.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_168.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_168.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_176.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_176.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_184.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_184.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_192.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_192.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_200.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_200.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_208.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_208.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_216.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_216.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_224.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_224.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_232.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_232.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_240.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_240.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_248.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_248.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_256.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_256.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_264.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_264.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_272.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_272.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_280.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_280.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_288.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_288.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_296.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_296.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_304.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_304.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_312.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_312.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_320.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_320.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_328.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_328.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_336.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_336.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_344.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_344.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_352.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_352.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_360.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_360.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_368.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_368.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_376.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_376.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_384.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_384.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_73.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_73.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_153.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_153.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_161.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_161.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_169.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_169.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_177.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_177.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_185.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_185.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_193.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_193.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_201.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_201.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_209.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_209.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_217.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_217.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_225.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_225.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_233.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_233.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_241.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_241.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_249.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_249.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_257.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_257.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_265.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_265.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_273.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_273.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_281.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_281.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_289.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_289.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_297.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_297.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_305.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_305.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_313.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_313.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_321.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_321.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_329.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_329.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_337.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_337.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_345.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_345.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_353.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_353.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_377.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_377.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_385.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_385.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_21.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_27.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_27.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_35.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_35.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_53.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_53.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_67.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_67.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_69.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_69.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_83.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_83.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_85.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_85.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_99.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_99.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_101.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_101.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_103.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_103.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_107.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_107.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_139.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_139.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_147.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_147.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_149.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_149.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_151.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_151.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_153.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_153.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_155.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_155.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_157.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_157.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_159.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_159.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_161.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_161.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_163.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_163.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_165.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_165.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_167.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_167.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_169.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_169.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_171.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_171.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_173.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_173.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_175.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_175.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_177.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_177.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_179.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_179.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_181.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_181.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_183.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_183.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_185.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_185.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_187.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_187.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_189.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_189.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_191.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_191.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_193.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_193.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_195.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_195.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_197.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_197.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_199.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_199.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_201.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_201.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_203.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_203.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_205.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_205.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_207.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_207.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_209.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_209.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_211.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_211.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_213.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_213.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_215.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_215.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_217.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_217.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_219.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_219.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_221.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_221.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_223.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_223.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_225.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_225.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_227.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_227.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_229.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_229.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_231.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_231.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_233.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_233.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_235.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_235.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_237.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_237.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_239.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_239.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_241.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_241.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_243.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_243.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_245.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_245.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_247.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_247.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_249.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_249.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_251.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_251.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_253.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_253.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_255.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_255.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_257.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_257.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_259.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_259.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_261.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_261.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_263.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_263.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_265.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_265.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_267.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_267.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_269.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_269.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_271.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_271.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_273.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_273.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_275.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_275.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_277.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_277.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_279.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_279.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_281.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_281.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_283.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_283.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_285.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_285.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_287.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_287.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_289.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_289.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_291.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_291.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_293.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_293.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_295.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_295.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_297.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_297.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_299.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_299.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_301.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_301.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_303.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_303.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_305.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_305.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_307.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_307.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_309.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_309.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_311.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_311.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_313.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_313.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_315.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_315.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_317.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_317.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_319.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_319.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_321.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_321.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_323.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_323.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_325.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_325.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_327.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_327.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_329.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_329.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_331.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_331.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_333.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_333.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_335.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_335.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_337.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_337.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_339.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_339.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_341.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_341.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_343.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_343.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_345.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_345.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_347.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_347.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_349.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_349.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_351.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_351.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_353.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_353.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_355.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_355.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_357.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_357.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_359.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_359.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_361.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_361.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_363.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_363.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_365.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_365.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_367.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_367.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_369.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_369.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_371.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_371.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_373.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_373.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_375.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_375.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_377.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_377.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_379.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_379.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_381.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_381.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_383.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_383.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_385.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_385.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_217.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_217.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_235.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_235.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_253.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_253.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_271.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_271.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_289.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_289.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_307.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_307.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_325.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_325.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_343.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_343.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_379.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_379.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_147.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_147.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_149.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_149.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_151.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_151.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_153.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_153.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_155.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_155.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_157.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_157.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_159.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_159.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_163.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_163.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_165.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_165.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_167.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_167.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_169.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_169.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_171.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_171.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_173.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_173.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_175.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_175.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_177.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_177.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_181.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_181.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_183.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_183.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_185.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_185.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_187.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_187.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_189.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_189.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_191.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_191.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_193.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_193.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_195.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_195.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_197.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_197.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_199.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_199.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_201.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_201.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_203.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_203.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_205.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_205.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_207.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_207.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_209.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_209.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_211.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_211.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_213.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_213.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_217.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_217.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_219.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_219.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_221.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_221.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_223.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_223.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_225.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_225.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_227.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_227.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_229.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_229.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_231.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_231.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_235.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_235.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_237.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_237.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_239.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_239.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_241.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_241.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_243.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_243.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_245.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_245.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_247.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_247.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_249.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_249.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_253.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_253.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_255.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_255.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_257.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_257.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_259.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_259.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_261.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_261.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_263.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_263.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_265.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_265.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_267.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_267.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_271.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_271.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_273.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_273.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_275.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_275.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_277.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_277.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_279.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_279.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_281.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_281.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_283.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_283.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_285.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_285.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_289.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_289.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_291.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_291.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_293.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_293.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_295.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_295.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_297.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_297.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_299.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_299.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_301.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_301.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_303.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_303.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_307.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_307.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_309.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_309.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_311.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_311.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_313.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_313.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_315.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_315.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_317.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_317.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_319.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_319.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_321.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_321.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_325.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_325.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_327.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_327.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_329.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_329.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_331.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_331.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_333.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_333.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_335.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_335.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_337.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_337.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_339.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_339.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_343.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_343.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_345.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_345.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_347.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_347.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_349.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_349.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_351.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_351.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_353.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_353.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_355.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_355.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_357.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_357.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_361.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_361.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_363.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_363.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_365.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_365.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_367.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_367.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_369.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_369.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_371.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_371.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_373.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_373.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_375.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_375.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_377.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_377.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_379.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_379.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_381.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_381.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_383.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_383.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_385.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_385.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:6] = 7'b0101110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:6] = 7'b1010001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:6] = 7'b0111111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:6] = 7'b1000000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:6] = 7'b0110100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:6] = 7'b1001011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_89.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_89.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_89.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_89.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:6] = 7'b0100111;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:6] = 7'b1011000;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_out[0:6] = 7'b0101101;
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_outb[0:6] = 7'b1010010;
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_out[0:6] = 7'b0001001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_outb[0:6] = 7'b1110110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_out[0:6] = 7'b0000111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_outb[0:6] = 7'b1111000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_out[0:6] = 7'b0101111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_outb[0:6] = 7'b1010000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_out[0:6] = 7'b0001010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_outb[0:6] = 7'b1110101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_8.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_8.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_9.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_9.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_10.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_10.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_11.mem_out[0:6] = 7'b0101010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_11.mem_outb[0:6] = 7'b1010101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_12.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_12.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_13.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_13.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_14.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_14.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_15.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_15.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_16.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_16.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_17.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_17.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_18.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_18.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_19.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_19.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_20.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_20.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_21.mem_out[0:6] = 7'b0110101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_21.mem_outb[0:6] = 7'b1001010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_22.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_22.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_23.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_23.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_24.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_24.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_25.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_25.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_26.mem_out[0:6] = 7'b0000110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_26.mem_outb[0:6] = 7'b1111001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_27.mem_out[0:6] = 7'b0111001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_27.mem_outb[0:6] = 7'b1000110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_28.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_28.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_29.mem_out[0:6] = 7'b0100111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_29.mem_outb[0:6] = 7'b1011000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_30.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_30.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_31.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_31.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_32.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_32.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_33.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_33.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_34.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_34.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_35.mem_out[0:6] = 7'b0000111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_35.mem_outb[0:6] = 7'b1111000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_36.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_36.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_37.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_37.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_38.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_38.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_39.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_39.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_40.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_40.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_41.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_41.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_42.mem_out[0:6] = 7'b0001010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_42.mem_outb[0:6] = 7'b1110101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_43.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_43.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_44.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_44.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_45.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_45.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_46.mem_out[0:6] = 7'b0110000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_46.mem_outb[0:6] = 7'b1001111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_47.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_47.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_48.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_48.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_49.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_49.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_50.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_50.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_51.mem_out[0:6] = 7'b0110001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_51.mem_outb[0:6] = 7'b1001110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_52.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_52.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_53.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_53.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_54.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_54.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_55.mem_out[0:6] = 7'b0000111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_55.mem_outb[0:6] = 7'b1111000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_56.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_56.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_57.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_57.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_58.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_58.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_59.mem_out[0:6] = 7'b0101000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_59.mem_outb[0:6] = 7'b1010111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_60.mem_out[0:6] = 7'b0011101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_60.mem_outb[0:6] = 7'b1100010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_61.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_61.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_62.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_62.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_63.mem_out[0:6] = 7'b0101110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_63.mem_outb[0:6] = 7'b1010001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_64.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_64.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_65.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_65.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_66.mem_out[0:6] = 7'b0110000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_66.mem_outb[0:6] = 7'b1001111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_67.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_67.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_68.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_68.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_69.mem_out[0:6] = 7'b0111100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_69.mem_outb[0:6] = 7'b1000011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_70.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_70.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_71.mem_out[0:6] = 7'b0101001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_71.mem_outb[0:6] = 7'b1010110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_72.mem_out[0:6] = 7'b0000110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_72.mem_outb[0:6] = 7'b1111001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_73.mem_out[0:6] = 7'b0011011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_73.mem_outb[0:6] = 7'b1100100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_74.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_74.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_75.mem_out[0:6] = 7'b0111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_75.mem_outb[0:6] = 7'b1000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_76.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_76.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_77.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_77.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_78.mem_out[0:6] = 7'b0001001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_78.mem_outb[0:6] = 7'b1110110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_79.mem_out[0:6] = 7'b0110101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_79.mem_outb[0:6] = 7'b1001010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_80.mem_out[0:6] = 7'b0001010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_80.mem_outb[0:6] = 7'b1110101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_81.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_81.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_82.mem_out[0:6] = 7'b0111101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_82.mem_outb[0:6] = 7'b1000010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_83.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_83.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_84.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_84.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_85.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_85.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_86.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_86.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_87.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_87.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_88.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_88.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_out[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_outb[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_out[0:6] = 7'b0011101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_outb[0:6] = 7'b1100010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_10.mem_out[0:6] = 7'b0000110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_10.mem_outb[0:6] = 7'b1111001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_11.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_11.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_12.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_12.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_13.mem_out[0:6] = 7'b0011011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_13.mem_outb[0:6] = 7'b1100100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_14.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_14.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_15.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_15.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_16.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_16.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_17.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_17.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_18.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_18.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_19.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_19.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_20.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_20.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_21.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_21.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_22.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_22.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_23.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_23.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_24.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_24.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_25.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_25.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_26.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_26.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_27.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_27.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_28.mem_out[0:6] = 7'b0011101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_28.mem_outb[0:6] = 7'b1100010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_29.mem_out[0:6] = 7'b0001010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_29.mem_outb[0:6] = 7'b1110101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_30.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_30.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_31.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_31.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_32.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_32.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_33.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_33.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_34.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_34.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_35.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_35.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_36.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_36.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_37.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_37.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_38.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_38.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_39.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_39.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_40.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_40.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_41.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_41.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_42.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_42.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_43.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_43.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_44.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_44.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_45.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_45.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_46.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_46.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_47.mem_out[0:6] = 7'b0000110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_47.mem_outb[0:6] = 7'b1111001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_48.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_48.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_49.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_49.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_50.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_50.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_51.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_51.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_52.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_52.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_53.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_53.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_54.mem_out[0:6] = 7'b0110001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_54.mem_outb[0:6] = 7'b1001110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_55.mem_out[0:6] = 7'b0101001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_55.mem_outb[0:6] = 7'b1010110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_56.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_56.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_57.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_57.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_58.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_58.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_59.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_59.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_60.mem_out[0:6] = 7'b0010000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_60.mem_outb[0:6] = 7'b1101111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_61.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_61.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_62.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_62.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_63.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_63.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_64.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_64.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_65.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_65.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_66.mem_out[0:6] = 7'b0111010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_66.mem_outb[0:6] = 7'b1000101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_67.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_67.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_68.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_68.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_69.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_69.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_70.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_70.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_71.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_71.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_72.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_72.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_73.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_73.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_74.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_74.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_75.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_75.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_76.mem_out[0:6] = 7'b0011011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_76.mem_outb[0:6] = 7'b1100100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_77.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_77.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_78.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_78.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_79.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_79.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_80.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_80.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_81.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_81.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_82.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_82.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_83.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_83.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_84.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_84.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_85.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_85.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_86.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_86.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_87.mem_out[0:6] = 7'b0000111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_87.mem_outb[0:6] = 7'b1111000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_88.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_88.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_89.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_89.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_89.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_89.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:6] = 7'b0100001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:6] = 7'b1011110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_out[0:6] = 7'b0001010;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_outb[0:6] = 7'b1110101;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:6] = 7'b0110010;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:6] = 7'b1001101;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:6] = 7'b0101110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:6] = 7'b1010001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:6] = 7'b0110000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:6] = 7'b1001111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:6] = 7'b0111000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:6] = 7'b1000111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_out[0:6] = 7'b0010000;
	force U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_outb[0:6] = 7'b1101111;
	force U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:6] = 7'b0101011;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:6] = 7'b1010100;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_out[0:6] = 7'b0101011;
	force U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_outb[0:6] = 7'b1010100;
	force U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_out[0:6] = 7'b0100010;
	force U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_outb[0:6] = 7'b1011101;
	force U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cby_2__4_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_out[0:6] = 7'b0110001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_outb[0:6] = 7'b1001110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_out[0:6] = 7'b0101001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_outb[0:6] = 7'b1010110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_out[0:6] = 7'b0010000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_outb[0:6] = 7'b1101111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_out[0:6] = 7'b0010000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_outb[0:6] = 7'b1101111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_8.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_8.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_9.mem_out[0:6] = 7'b0101000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_9.mem_outb[0:6] = 7'b1010111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_10.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_10.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_11.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_11.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_12.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_12.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_13.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_13.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_14.mem_out[0:6] = 7'b0010000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_14.mem_outb[0:6] = 7'b1101111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_15.mem_out[0:6] = 7'b0100000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_15.mem_outb[0:6] = 7'b1011111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_16.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_16.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_17.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_17.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_18.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_18.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_19.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_19.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_20.mem_out[0:6] = 7'b0100000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_20.mem_outb[0:6] = 7'b1011111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_21.mem_out[0:6] = 7'b0100111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_21.mem_outb[0:6] = 7'b1011000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_22.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_22.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_23.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_23.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_24.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_24.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_25.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_25.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_26.mem_out[0:6] = 7'b0111000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_26.mem_outb[0:6] = 7'b1000111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_27.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_27.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_28.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_28.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_29.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_29.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_30.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_30.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_31.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_31.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_32.mem_out[0:6] = 7'b0011101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_32.mem_outb[0:6] = 7'b1100010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_33.mem_out[0:6] = 7'b0000111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_33.mem_outb[0:6] = 7'b1111000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_34.mem_out[0:6] = 7'b0000110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_34.mem_outb[0:6] = 7'b1111001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_35.mem_out[0:6] = 7'b0010111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_35.mem_outb[0:6] = 7'b1101000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_36.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_36.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_37.mem_out[0:6] = 7'b0011011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_37.mem_outb[0:6] = 7'b1100100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_38.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_38.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_39.mem_out[0:6] = 7'b0101101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_39.mem_outb[0:6] = 7'b1010010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_40.mem_out[0:6] = 7'b0001001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_40.mem_outb[0:6] = 7'b1110110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_41.mem_out[0:6] = 7'b0011011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_41.mem_outb[0:6] = 7'b1100100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_42.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_42.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_43.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_43.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_44.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_44.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_45.mem_out[0:6] = 7'b0100111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_45.mem_outb[0:6] = 7'b1011000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_46.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_46.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_47.mem_out[0:6] = 7'b0110101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_47.mem_outb[0:6] = 7'b1001010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_48.mem_out[0:6] = 7'b0100111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_48.mem_outb[0:6] = 7'b1011000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_49.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_49.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_50.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_50.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_51.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_51.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_52.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_52.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_53.mem_out[0:6] = 7'b0111001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_53.mem_outb[0:6] = 7'b1000110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_54.mem_out[0:6] = 7'b0110000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_54.mem_outb[0:6] = 7'b1001111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_55.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_55.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_56.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_56.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_57.mem_out[0:6] = 7'b0101011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_57.mem_outb[0:6] = 7'b1010100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_58.mem_out[0:6] = 7'b0101101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_58.mem_outb[0:6] = 7'b1010010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_59.mem_out[0:6] = 7'b0100011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_59.mem_outb[0:6] = 7'b1011100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_60.mem_out[0:6] = 7'b0100110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_60.mem_outb[0:6] = 7'b1011001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_61.mem_out[0:6] = 7'b0000110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_61.mem_outb[0:6] = 7'b1111001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_62.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_62.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_63.mem_out[0:6] = 7'b0111111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_63.mem_outb[0:6] = 7'b1000000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_64.mem_out[0:6] = 7'b0011110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_64.mem_outb[0:6] = 7'b1100001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_65.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_65.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_66.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_66.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_67.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_67.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_68.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_68.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_69.mem_out[0:6] = 7'b0110110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_69.mem_outb[0:6] = 7'b1001001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_70.mem_out[0:6] = 7'b0111000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_70.mem_outb[0:6] = 7'b1000111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_71.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_71.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_72.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_72.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_73.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_73.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_74.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_74.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_75.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_75.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_76.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_76.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_77.mem_out[0:6] = 7'b0010011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_77.mem_outb[0:6] = 7'b1101100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_78.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_78.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_79.mem_out[0:6] = 7'b0011101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_79.mem_outb[0:6] = 7'b1100010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_80.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_80.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_81.mem_out[0:6] = 7'b0100101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_81.mem_outb[0:6] = 7'b1011010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_82.mem_out[0:6] = 7'b0111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_82.mem_outb[0:6] = 7'b1000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_83.mem_out[0:6] = 7'b0011101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_83.mem_outb[0:6] = 7'b1100010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_84.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_84.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_85.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_85.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_86.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_86.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_87.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_87.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_88.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_88.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_out[0:6] = 7'b0100110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_outb[0:6] = 7'b1011001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_out[0:6] = 7'b0100101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_outb[0:6] = 7'b1011010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_out[0:6] = 7'b0110100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_outb[0:6] = 7'b1001011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_out[0:6] = 7'b0100001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_outb[0:6] = 7'b1011110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_out[0:6] = 7'b0000111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_outb[0:6] = 7'b1111000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_out[0:6] = 7'b0001111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_outb[0:6] = 7'b1110000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_out[0:6] = 7'b0001010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_outb[0:6] = 7'b1110101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_10.mem_out[0:6] = 7'b0100000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_10.mem_outb[0:6] = 7'b1011111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_11.mem_out[0:6] = 7'b0000100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_11.mem_outb[0:6] = 7'b1111011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_12.mem_out[0:6] = 7'b0101010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_12.mem_outb[0:6] = 7'b1010101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_13.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_13.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_14.mem_out[0:6] = 7'b0110101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_14.mem_outb[0:6] = 7'b1001010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_15.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_15.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_16.mem_out[0:6] = 7'b0100010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_16.mem_outb[0:6] = 7'b1011101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_17.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_17.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_18.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_18.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_19.mem_out[0:6] = 7'b0011100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_19.mem_outb[0:6] = 7'b1100011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_20.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_20.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_21.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_21.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_22.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_22.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_23.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_23.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_24.mem_out[0:6] = 7'b0010010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_24.mem_outb[0:6] = 7'b1101101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_25.mem_out[0:6] = 7'b0010001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_25.mem_outb[0:6] = 7'b1101110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_26.mem_out[0:6] = 7'b0110110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_26.mem_outb[0:6] = 7'b1001001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_27.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_27.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_28.mem_out[0:6] = 7'b1101111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_28.mem_outb[0:6] = 7'b0010000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_29.mem_out[0:6] = 7'b0101111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_29.mem_outb[0:6] = 7'b1010000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_30.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_30.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_31.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_31.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_32.mem_out[0:6] = 7'b0110011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_32.mem_outb[0:6] = 7'b1001100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_33.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_33.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_34.mem_out[0:6] = 7'b0000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_34.mem_outb[0:6] = 7'b1111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_35.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_35.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_36.mem_out[0:6] = 7'b0101101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_36.mem_outb[0:6] = 7'b1010010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_37.mem_out[0:6] = 7'b0110011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_37.mem_outb[0:6] = 7'b1001100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_38.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_38.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_39.mem_out[0:6] = 7'b0111111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_39.mem_outb[0:6] = 7'b1000000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_40.mem_out[0:6] = 7'b0100101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_40.mem_outb[0:6] = 7'b1011010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_41.mem_out[0:6] = 7'b0011011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_41.mem_outb[0:6] = 7'b1100100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_42.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_42.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_43.mem_out[0:6] = 7'b0110111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_43.mem_outb[0:6] = 7'b1001000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_44.mem_out[0:6] = 7'b0110001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_44.mem_outb[0:6] = 7'b1001110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_45.mem_out[0:6] = 7'b0001101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_45.mem_outb[0:6] = 7'b1110010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_46.mem_out[0:6] = 7'b0011011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_46.mem_outb[0:6] = 7'b1100100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_47.mem_out[0:6] = 7'b0100100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_47.mem_outb[0:6] = 7'b1011011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_48.mem_out[0:6] = 7'b0011101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_48.mem_outb[0:6] = 7'b1100010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_49.mem_out[0:6] = 7'b0010100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_49.mem_outb[0:6] = 7'b1101011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_50.mem_out[0:6] = 7'b0011001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_50.mem_outb[0:6] = 7'b1100110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_51.mem_out[0:6] = 7'b0100011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_51.mem_outb[0:6] = 7'b1011100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_52.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_52.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_53.mem_out[0:6] = 7'b0001100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_53.mem_outb[0:6] = 7'b1110011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_54.mem_out[0:6] = 7'b0001110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_54.mem_outb[0:6] = 7'b1110001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_55.mem_out[0:6] = 7'b0010000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_55.mem_outb[0:6] = 7'b1101111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_56.mem_out[0:6] = 7'b0110010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_56.mem_outb[0:6] = 7'b1001101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_57.mem_out[0:6] = 7'b0110011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_57.mem_outb[0:6] = 7'b1001100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_58.mem_out[0:6] = 7'b0010101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_58.mem_outb[0:6] = 7'b1101010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_59.mem_out[0:6] = 7'b0100011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_59.mem_outb[0:6] = 7'b1011100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_60.mem_out[0:6] = 7'b0101100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_60.mem_outb[0:6] = 7'b1010011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_61.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_61.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_62.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_62.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_63.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_63.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_64.mem_out[0:6] = 7'b0100100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_64.mem_outb[0:6] = 7'b1011011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_65.mem_out[0:6] = 7'b0000010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_65.mem_outb[0:6] = 7'b1111101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_66.mem_out[0:6] = 7'b0001010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_66.mem_outb[0:6] = 7'b1110101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_67.mem_out[0:6] = 7'b0101110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_67.mem_outb[0:6] = 7'b1010001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_68.mem_out[0:6] = 7'b0110000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_68.mem_outb[0:6] = 7'b1001111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_69.mem_out[0:6] = 7'b0000101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_69.mem_outb[0:6] = 7'b1111010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_70.mem_out[0:6] = 7'b0000110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_70.mem_outb[0:6] = 7'b1111001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_71.mem_out[0:6] = 7'b0101101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_71.mem_outb[0:6] = 7'b1010010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_72.mem_out[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_72.mem_outb[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_73.mem_out[0:6] = 7'b0001011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_73.mem_outb[0:6] = 7'b1110100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_74.mem_out[0:6] = 7'b1011111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_74.mem_outb[0:6] = 7'b0100000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_75.mem_out[0:6] = 7'b0111011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_75.mem_outb[0:6] = 7'b1000100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_76.mem_out[0:6] = 7'b0011000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_76.mem_outb[0:6] = 7'b1100111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_77.mem_out[0:6] = 7'b0111111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_77.mem_outb[0:6] = 7'b1000000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_78.mem_out[0:6] = 7'b0101110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_78.mem_outb[0:6] = 7'b1010001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_79.mem_out[0:6] = 7'b0011010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_79.mem_outb[0:6] = 7'b1100101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_80.mem_out[0:6] = 7'b0010110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_80.mem_outb[0:6] = 7'b1101001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_81.mem_out[0:6] = 7'b0101111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_81.mem_outb[0:6] = 7'b1010000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_82.mem_out[0:6] = 7'b0100110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_82.mem_outb[0:6] = 7'b1011001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_83.mem_out[0:6] = 7'b0001001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_83.mem_outb[0:6] = 7'b1110110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_84.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_84.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_85.mem_out[0:6] = 7'b0100001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_85.mem_outb[0:6] = 7'b1011110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_86.mem_out[0:6] = 7'b0111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_86.mem_outb[0:6] = 7'b1000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_87.mem_out[0:6] = 7'b0000011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_87.mem_outb[0:6] = 7'b1111100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_88.mem_out[0:6] = 7'b0001000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_88.mem_outb[0:6] = 7'b1110111;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_8.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_8.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_9.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_9.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_10.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_10.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_11.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_11.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_12.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_12.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_13.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_13.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_14.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_14.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_15.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_15.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_16.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_16.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_17.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_17.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_18.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_18.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_19.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_19.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_20.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_20.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_21.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_21.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_22.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_22.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_23.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_23.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_24.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_24.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_25.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_25.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_26.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_26.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_27.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_27.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_28.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_28.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_29.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_29.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_30.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_30.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_31.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_31.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_32.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_32.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_33.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_33.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_34.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_34.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_35.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_35.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_36.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_36.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_37.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_37.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_38.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_38.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_39.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_39.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_40.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_40.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_41.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_41.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_42.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_42.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_43.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_43.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_44.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_44.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_45.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_45.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_46.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_46.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_47.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_47.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_48.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_48.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_49.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_49.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_50.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_50.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_51.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_51.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_52.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_52.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_53.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_53.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_54.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_54.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_55.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_55.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_56.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_56.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_57.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_57.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_58.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_58.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_59.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_59.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_60.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_60.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_61.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_61.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_62.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_62.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_63.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_63.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_64.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_64.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_65.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_65.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_66.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_66.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_67.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_67.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_68.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_68.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_69.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_69.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_70.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_70.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_71.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_71.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_72.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_72.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_73.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_73.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_74.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_74.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_75.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_75.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_76.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_76.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_77.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_77.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_78.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_78.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_79.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_79.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_80.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_80.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_81.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_81.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_82.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_82.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_83.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_83.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_84.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_84.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_85.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_85.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_86.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_86.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_87.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_87.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_88.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_88.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_2.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_3.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_3.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_4.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_4.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_5.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_5.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_6.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_6.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_7.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_7.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_outb[0:6] = {7{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_out[0:6] = {7{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_outb[0:6] = {7{1'b1}};
end
// ----- End assign bitstream to configuration memories -----
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for router_tb_top_formal_verification -----

//----- Default net type -----
`default_nettype wire

