//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[10][3]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Jul 24 20:28:26 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_10__3_ -----
module sb_10__3_(prog_clk,
                 chany_top_in,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                 chany_bottom_in,
                 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                 chanx_left_in,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                 ccff_head,
                 chany_top_out,
                 chany_bottom_out,
                 chanx_left_out,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:104] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:104] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:104] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:104] chany_top_out;
//----- OUTPUT PORTS -----
output [0:104] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:104] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_16_sram;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_17_sram;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_18_sram;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_19_sram;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_20_sram;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_21_sram;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_22_sram;
wire [0:1] mux_tree_tapbuf_size2_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_23_sram;
wire [0:1] mux_tree_tapbuf_size2_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_24_sram;
wire [0:1] mux_tree_tapbuf_size2_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_25_sram;
wire [0:1] mux_tree_tapbuf_size2_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_26_sram;
wire [0:1] mux_tree_tapbuf_size2_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_27_sram;
wire [0:1] mux_tree_tapbuf_size2_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_28_sram;
wire [0:1] mux_tree_tapbuf_size2_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_29_sram;
wire [0:1] mux_tree_tapbuf_size2_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_30_sram;
wire [0:1] mux_tree_tapbuf_size2_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_31_sram;
wire [0:1] mux_tree_tapbuf_size2_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_32_sram;
wire [0:1] mux_tree_tapbuf_size2_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_33_sram;
wire [0:1] mux_tree_tapbuf_size2_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_34_sram;
wire [0:1] mux_tree_tapbuf_size2_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_35_sram;
wire [0:1] mux_tree_tapbuf_size2_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_36_sram;
wire [0:1] mux_tree_tapbuf_size2_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_37_sram;
wire [0:1] mux_tree_tapbuf_size2_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_38_sram;
wire [0:1] mux_tree_tapbuf_size2_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_39_sram;
wire [0:1] mux_tree_tapbuf_size2_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_40_sram;
wire [0:1] mux_tree_tapbuf_size2_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_41_sram;
wire [0:1] mux_tree_tapbuf_size2_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_42_sram;
wire [0:1] mux_tree_tapbuf_size2_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_43_sram;
wire [0:1] mux_tree_tapbuf_size2_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_44_sram;
wire [0:1] mux_tree_tapbuf_size2_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_45_sram;
wire [0:1] mux_tree_tapbuf_size2_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_46_sram;
wire [0:1] mux_tree_tapbuf_size2_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_47_sram;
wire [0:1] mux_tree_tapbuf_size2_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_48_sram;
wire [0:1] mux_tree_tapbuf_size2_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_49_sram;
wire [0:1] mux_tree_tapbuf_size2_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_50_sram;
wire [0:1] mux_tree_tapbuf_size2_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_51_sram;
wire [0:1] mux_tree_tapbuf_size2_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_52_sram;
wire [0:1] mux_tree_tapbuf_size2_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_53_sram;
wire [0:1] mux_tree_tapbuf_size2_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_54_sram;
wire [0:1] mux_tree_tapbuf_size2_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_55_sram;
wire [0:1] mux_tree_tapbuf_size2_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_56_sram;
wire [0:1] mux_tree_tapbuf_size2_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_57_sram;
wire [0:1] mux_tree_tapbuf_size2_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_58_sram;
wire [0:1] mux_tree_tapbuf_size2_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_59_sram;
wire [0:1] mux_tree_tapbuf_size2_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_60_sram;
wire [0:1] mux_tree_tapbuf_size2_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_61_sram;
wire [0:1] mux_tree_tapbuf_size2_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_62_sram;
wire [0:1] mux_tree_tapbuf_size2_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_63_sram;
wire [0:1] mux_tree_tapbuf_size2_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_64_sram;
wire [0:1] mux_tree_tapbuf_size2_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_65_sram;
wire [0:1] mux_tree_tapbuf_size2_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_66_sram;
wire [0:1] mux_tree_tapbuf_size2_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_67_sram;
wire [0:1] mux_tree_tapbuf_size2_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_68_sram;
wire [0:1] mux_tree_tapbuf_size2_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_69_sram;
wire [0:1] mux_tree_tapbuf_size2_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_70_sram;
wire [0:1] mux_tree_tapbuf_size2_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_71_sram;
wire [0:1] mux_tree_tapbuf_size2_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_72_sram;
wire [0:1] mux_tree_tapbuf_size2_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_73_sram;
wire [0:1] mux_tree_tapbuf_size2_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_74_sram;
wire [0:1] mux_tree_tapbuf_size2_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_75_sram;
wire [0:1] mux_tree_tapbuf_size2_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_76_sram;
wire [0:1] mux_tree_tapbuf_size2_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_77_sram;
wire [0:1] mux_tree_tapbuf_size2_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_78_sram;
wire [0:1] mux_tree_tapbuf_size2_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_79_sram;
wire [0:1] mux_tree_tapbuf_size2_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_80_sram;
wire [0:1] mux_tree_tapbuf_size2_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_81_sram;
wire [0:1] mux_tree_tapbuf_size2_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_82_sram;
wire [0:1] mux_tree_tapbuf_size2_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_4_sram;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_5_sram;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_6_sram;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_29_sram;
wire [0:2] mux_tree_tapbuf_size5_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_30_sram;
wire [0:2] mux_tree_tapbuf_size5_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_31_sram;
wire [0:2] mux_tree_tapbuf_size5_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_32_sram;
wire [0:2] mux_tree_tapbuf_size5_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_33_sram;
wire [0:2] mux_tree_tapbuf_size5_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_34_sram;
wire [0:2] mux_tree_tapbuf_size5_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_35_sram;
wire [0:2] mux_tree_tapbuf_size5_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_36_sram;
wire [0:2] mux_tree_tapbuf_size5_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_37_sram;
wire [0:2] mux_tree_tapbuf_size5_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_38_sram;
wire [0:2] mux_tree_tapbuf_size5_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_39_sram;
wire [0:2] mux_tree_tapbuf_size5_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_40_sram;
wire [0:2] mux_tree_tapbuf_size5_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_41_sram;
wire [0:2] mux_tree_tapbuf_size5_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_42_sram;
wire [0:2] mux_tree_tapbuf_size5_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_43_sram;
wire [0:2] mux_tree_tapbuf_size5_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_44_sram;
wire [0:2] mux_tree_tapbuf_size5_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_45_sram;
wire [0:2] mux_tree_tapbuf_size5_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_46_sram;
wire [0:2] mux_tree_tapbuf_size5_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_47_sram;
wire [0:2] mux_tree_tapbuf_size5_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size5 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[0], chanx_left_in[27], chanx_left_in[54], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size5 mux_top_track_32 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[23], chanx_left_in[50], chanx_left_in[77], chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size5 mux_top_track_40 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[22], chanx_left_in[49], chanx_left_in[76], chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size5 mux_top_track_48 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[21], chanx_left_in[48], chanx_left_in[75], chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size5 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[20], chanx_left_in[47], chanx_left_in[74], chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size5 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[19], chanx_left_in[46], chanx_left_in[73], chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size5 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[18], chanx_left_in[45], chanx_left_in[72], chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size5 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[17], chanx_left_in[44], chanx_left_in[71], chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size5 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[16], chanx_left_in[43], chanx_left_in[70], chanx_left_in[97]}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size5 mux_top_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[15], chanx_left_in[42], chanx_left_in[69], chanx_left_in[96]}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size5 mux_top_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[14], chanx_left_in[41], chanx_left_in[68], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size5 mux_top_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[13], chanx_left_in[40], chanx_left_in[67], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size5 mux_top_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[12], chanx_left_in[39], chanx_left_in[66], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size5 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[11], chanx_left_in[38], chanx_left_in[65], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size5 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[10], chanx_left_in[37], chanx_left_in[64], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size5 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[9], chanx_left_in[36], chanx_left_in[63], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size5 mux_top_track_152 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[8], chanx_left_in[35], chanx_left_in[62], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size5 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[7], chanx_left_in[34], chanx_left_in[61], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size5 mux_top_track_168 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[6], chanx_left_in[33], chanx_left_in[60], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size5 mux_top_track_176 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[5], chanx_left_in[32], chanx_left_in[59], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size5 mux_top_track_184 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[4], chanx_left_in[31], chanx_left_in[58], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size5 mux_top_track_192 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[3], chanx_left_in[30], chanx_left_in[57], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size5 mux_top_track_200 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[2], chanx_left_in[29], chanx_left_in[56], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size5 mux_top_track_208 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[1], chanx_left_in[28], chanx_left_in[55], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size5 mux_bottom_track_1 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[1], chanx_left_in[28], chanx_left_in[55], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size5 mux_bottom_track_9 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[2], chanx_left_in[29], chanx_left_in[56], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size5 mux_bottom_track_17 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[3], chanx_left_in[30], chanx_left_in[57], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size5 mux_bottom_track_25 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[4], chanx_left_in[31], chanx_left_in[58], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size5 mux_bottom_track_33 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[5], chanx_left_in[32], chanx_left_in[59], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size5 mux_bottom_track_41 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[6], chanx_left_in[33], chanx_left_in[60], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_size5_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_29_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size5 mux_bottom_track_49 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[7], chanx_left_in[34], chanx_left_in[61], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_size5_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_30_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size5 mux_bottom_track_57 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[8], chanx_left_in[35], chanx_left_in[62], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_size5_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_31_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size5 mux_bottom_track_65 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[9], chanx_left_in[36], chanx_left_in[63], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_size5_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_32_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size5 mux_bottom_track_73 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[10], chanx_left_in[37], chanx_left_in[64], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_size5_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_33_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size5 mux_bottom_track_81 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[11], chanx_left_in[38], chanx_left_in[65], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_size5_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_34_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size5 mux_bottom_track_89 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[12], chanx_left_in[39], chanx_left_in[66], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_size5_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_35_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size5 mux_bottom_track_97 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[13], chanx_left_in[40], chanx_left_in[67], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_size5_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_36_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size5 mux_bottom_track_105 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[14], chanx_left_in[41], chanx_left_in[68], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_size5_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_37_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size5 mux_bottom_track_113 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[15], chanx_left_in[42], chanx_left_in[69], chanx_left_in[96]}),
		.sram(mux_tree_tapbuf_size5_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_38_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size5 mux_bottom_track_121 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[16], chanx_left_in[43], chanx_left_in[70], chanx_left_in[97]}),
		.sram(mux_tree_tapbuf_size5_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_39_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size5 mux_bottom_track_129 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[17], chanx_left_in[44], chanx_left_in[71], chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size5_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_40_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size5 mux_bottom_track_137 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[18], chanx_left_in[45], chanx_left_in[72], chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size5_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_41_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size5 mux_bottom_track_145 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[19], chanx_left_in[46], chanx_left_in[73], chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size5_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_42_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size5 mux_bottom_track_153 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[20], chanx_left_in[47], chanx_left_in[74], chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size5_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_43_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size5 mux_bottom_track_161 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[21], chanx_left_in[48], chanx_left_in[75], chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size5_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_44_sram_inv[0:2]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size5 mux_bottom_track_169 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[22], chanx_left_in[49], chanx_left_in[76], chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size5_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_45_sram_inv[0:2]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size5 mux_bottom_track_177 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[23], chanx_left_in[50], chanx_left_in[77], chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size5_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_46_sram_inv[0:2]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size5 mux_bottom_track_209 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[0], chanx_left_in[27], chanx_left_in[54], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_size5_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_47_sram_inv[0:2]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size5_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_29_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_30_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_31_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_32_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_33_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_34_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_35_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_36_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_37_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_38_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_39_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_40_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_41_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_42_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_43_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_44_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_45_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_46_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_47_sram_inv[0:2]));

	mux_tree_tapbuf_size4 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[26], chanx_left_in[53], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size4 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[25], chanx_left_in[52], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size4 mux_top_track_24 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[24], chanx_left_in[51], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size4 mux_bottom_track_185 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[24], chanx_left_in[51], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size4 mux_bottom_track_193 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[25], chanx_left_in[52], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_size4_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_4_sram_inv[0:2]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size4 mux_bottom_track_201 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[26], chanx_left_in[53], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_size4_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_5_sram_inv[0:2]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size4 mux_left_track_163 (
		.in({chany_top_in[32], chany_top_in[99], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size4_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_6_sram_inv[0:2]),
		.out(chanx_left_out[81]));

	mux_tree_tapbuf_size4_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_4_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_5_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_163 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_6_sram_inv[0:2]));

	mux_tree_tapbuf_size3 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size3 mux_left_track_3 (
		.in({chany_bottom_in[0], chany_bottom_in[3], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_size3 mux_left_track_19 (
		.in({chany_bottom_in[10], chany_bottom_in[35], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_size3 mux_left_track_23 (
		.in({chany_bottom_in[13], chany_bottom_in[43], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_size3 mux_left_track_37 (
		.in({chany_bottom_in[22], chany_bottom_in[71], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_size3 mux_left_track_43 (
		.in({chany_bottom_in[26], chany_bottom_in[83], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_size3 mux_left_track_55 (
		.in({chany_bottom_in[34], chany_bottom_in[104], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_size3 mux_left_track_63 (
		.in({chany_top_in[98], chany_bottom_in[40], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_size3 mux_left_track_73 (
		.in({chany_top_in[92], chany_bottom_in[46], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size3 mux_left_track_83 (
		.in({chany_top_in[85], chany_bottom_in[53], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_size3 mux_left_track_91 (
		.in({chany_top_in[80], chany_bottom_in[58], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_size3 mux_left_track_103 (
		.in({chany_top_in[72], chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_size3 mux_left_track_109 (
		.in({chany_top_in[68], chany_bottom_in[70], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_size3 mux_left_track_123 (
		.in({chany_top_in[58], chany_bottom_in[80], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_size3 mux_left_track_127 (
		.in({chany_top_in[56], chany_bottom_in[82], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_size3 mux_left_track_143 (
		.in({chany_top_in[45], chany_bottom_in[93], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_size3 mux_left_track_145 (
		.in({chany_top_in[44], chany_bottom_in[94], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size3 mux_left_track_181 (
		.in({chany_top_in[20], chany_top_in[63], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chanx_left_out[90]));

	mux_tree_tapbuf_size3 mux_left_track_183 (
		.in({chany_top_in[18], chany_top_in[59], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_size3 mux_left_track_199 (
		.in({chany_top_in[8], chany_top_in[27], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chanx_left_out[99]));

	mux_tree_tapbuf_size3 mux_left_track_203 (
		.in({chany_top_in[5], chany_top_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chanx_left_out[101]));

	mux_tree_tapbuf_size3_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_181 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_183 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_199 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_203 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2 mux_left_track_5 (
		.in({chany_bottom_in[1], chany_bottom_in[7]}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_size2 mux_left_track_7 (
		.in({chany_bottom_in[2], chany_bottom_in[11]}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_size2 mux_left_track_9 (
		.in({chany_bottom_in[4], chany_bottom_in[15]}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size2 mux_left_track_11 (
		.in({chany_bottom_in[5], chany_bottom_in[19]}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_size2 mux_left_track_13 (
		.in({chany_bottom_in[6], chany_bottom_in[23]}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_size2 mux_left_track_15 (
		.in({chany_bottom_in[8], chany_bottom_in[27]}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_size2 mux_left_track_17 (
		.in({chany_bottom_in[9], chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size2 mux_left_track_21 (
		.in({chany_bottom_in[12], chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_size2 mux_left_track_25 (
		.in({chany_bottom_in[14], chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size2 mux_left_track_27 (
		.in({chany_bottom_in[16], chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_size2 mux_left_track_29 (
		.in({chany_bottom_in[17], chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_size2 mux_left_track_31 (
		.in({chany_bottom_in[18], chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_size2 mux_left_track_33 (
		.in({chany_bottom_in[20], chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size2 mux_left_track_35 (
		.in({chany_bottom_in[21], chany_bottom_in[67]}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_size2 mux_left_track_39 (
		.in({chany_bottom_in[24], chany_bottom_in[75]}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_size2 mux_left_track_41 (
		.in({chany_bottom_in[25], chany_bottom_in[79]}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size2 mux_left_track_45 (
		.in({chany_bottom_in[28], chany_bottom_in[87]}),
		.sram(mux_tree_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_16_sram_inv[0:1]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_size2 mux_left_track_47 (
		.in({chany_bottom_in[29], chany_bottom_in[91]}),
		.sram(mux_tree_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_17_sram_inv[0:1]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_size2 mux_left_track_49 (
		.in({chany_bottom_in[30], chany_bottom_in[95]}),
		.sram(mux_tree_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_18_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size2 mux_left_track_51 (
		.in({chany_bottom_in[32], chany_bottom_in[99]}),
		.sram(mux_tree_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_19_sram_inv[0:1]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_size2 mux_left_track_53 (
		.in({chany_bottom_in[33], chany_bottom_in[103]}),
		.sram(mux_tree_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_20_sram_inv[0:1]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_size2 mux_left_track_57 (
		.in({chany_top_in[102], chany_bottom_in[36]}),
		.sram(mux_tree_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_21_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size2 mux_left_track_59 (
		.in({chany_top_in[101], chany_bottom_in[37]}),
		.sram(mux_tree_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_22_sram_inv[0:1]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_size2 mux_left_track_61 (
		.in({chany_top_in[100], chany_bottom_in[38]}),
		.sram(mux_tree_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_23_sram_inv[0:1]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_size2 mux_left_track_65 (
		.in({chany_top_in[97], chany_bottom_in[41]}),
		.sram(mux_tree_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_24_sram_inv[0:1]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size2 mux_left_track_67 (
		.in({chany_top_in[96], chany_bottom_in[42]}),
		.sram(mux_tree_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_25_sram_inv[0:1]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_size2 mux_left_track_69 (
		.in({chany_top_in[94], chany_bottom_in[44]}),
		.sram(mux_tree_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_26_sram_inv[0:1]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_size2 mux_left_track_71 (
		.in({chany_top_in[93], chany_bottom_in[45]}),
		.sram(mux_tree_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_27_sram_inv[0:1]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_size2 mux_left_track_75 (
		.in({chany_top_in[90], chany_bottom_in[48]}),
		.sram(mux_tree_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_28_sram_inv[0:1]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_size2 mux_left_track_77 (
		.in({chany_top_in[89], chany_bottom_in[49]}),
		.sram(mux_tree_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_29_sram_inv[0:1]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_size2 mux_left_track_79 (
		.in({chany_top_in[88], chany_bottom_in[50]}),
		.sram(mux_tree_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_30_sram_inv[0:1]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_size2 mux_left_track_81 (
		.in({chany_top_in[86], chany_bottom_in[52]}),
		.sram(mux_tree_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_31_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size2 mux_left_track_85 (
		.in({chany_top_in[84], chany_bottom_in[54]}),
		.sram(mux_tree_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_32_sram_inv[0:1]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_size2 mux_left_track_87 (
		.in({chany_top_in[82], chany_bottom_in[56]}),
		.sram(mux_tree_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_33_sram_inv[0:1]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_size2 mux_left_track_89 (
		.in({chany_top_in[81], chany_bottom_in[57]}),
		.sram(mux_tree_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_34_sram_inv[0:1]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size2 mux_left_track_93 (
		.in({chany_top_in[78], chany_bottom_in[60]}),
		.sram(mux_tree_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_35_sram_inv[0:1]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_size2 mux_left_track_95 (
		.in({chany_top_in[77], chany_bottom_in[61]}),
		.sram(mux_tree_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_36_sram_inv[0:1]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_size2 mux_left_track_97 (
		.in({chany_top_in[76], chany_bottom_in[62]}),
		.sram(mux_tree_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_37_sram_inv[0:1]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size2 mux_left_track_99 (
		.in({chany_top_in[74], chany_bottom_in[64]}),
		.sram(mux_tree_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_38_sram_inv[0:1]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_size2 mux_left_track_101 (
		.in({chany_top_in[73], chany_bottom_in[65]}),
		.sram(mux_tree_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_39_sram_inv[0:1]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_size2 mux_left_track_105 (
		.in({chany_top_in[70], chany_bottom_in[68]}),
		.sram(mux_tree_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_40_sram_inv[0:1]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size2 mux_left_track_107 (
		.in({chany_top_in[69], chany_bottom_in[69]}),
		.sram(mux_tree_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_41_sram_inv[0:1]),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_size2 mux_left_track_111 (
		.in({chany_top_in[66], chany_bottom_in[72]}),
		.sram(mux_tree_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_42_sram_inv[0:1]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_size2 mux_left_track_113 (
		.in({chany_top_in[65], chany_bottom_in[73]}),
		.sram(mux_tree_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_43_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size2 mux_left_track_115 (
		.in({chany_top_in[64], chany_bottom_in[74]}),
		.sram(mux_tree_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_44_sram_inv[0:1]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_size2 mux_left_track_117 (
		.in({chany_top_in[62], chany_bottom_in[76]}),
		.sram(mux_tree_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_45_sram_inv[0:1]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_size2 mux_left_track_119 (
		.in({chany_top_in[61], chany_bottom_in[77]}),
		.sram(mux_tree_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_46_sram_inv[0:1]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_size2 mux_left_track_121 (
		.in({chany_top_in[60], chany_bottom_in[78]}),
		.sram(mux_tree_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_47_sram_inv[0:1]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size2 mux_left_track_125 (
		.in({chany_top_in[57], chany_bottom_in[81]}),
		.sram(mux_tree_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_48_sram_inv[0:1]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_size2 mux_left_track_129 (
		.in({chany_top_in[54], chany_bottom_in[84]}),
		.sram(mux_tree_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_49_sram_inv[0:1]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size2 mux_left_track_131 (
		.in({chany_top_in[53], chany_bottom_in[85]}),
		.sram(mux_tree_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_50_sram_inv[0:1]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_size2 mux_left_track_133 (
		.in({chany_top_in[52], chany_bottom_in[86]}),
		.sram(mux_tree_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_51_sram_inv[0:1]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_size2 mux_left_track_135 (
		.in({chany_top_in[50], chany_bottom_in[88]}),
		.sram(mux_tree_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_52_sram_inv[0:1]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_size2 mux_left_track_137 (
		.in({chany_top_in[49], chany_bottom_in[89]}),
		.sram(mux_tree_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_53_sram_inv[0:1]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size2 mux_left_track_139 (
		.in({chany_top_in[48], chany_bottom_in[90]}),
		.sram(mux_tree_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_54_sram_inv[0:1]),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_size2 mux_left_track_141 (
		.in({chany_top_in[46], chany_bottom_in[92]}),
		.sram(mux_tree_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_55_sram_inv[0:1]),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_size2 mux_left_track_147 (
		.in({chany_top_in[42], chany_bottom_in[96]}),
		.sram(mux_tree_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_56_sram_inv[0:1]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_size2 mux_left_track_149 (
		.in({chany_top_in[41], chany_bottom_in[97]}),
		.sram(mux_tree_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_57_sram_inv[0:1]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_size2 mux_left_track_151 (
		.in({chany_top_in[40], chany_bottom_in[98]}),
		.sram(mux_tree_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_58_sram_inv[0:1]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_size2 mux_left_track_153 (
		.in({chany_top_in[38], chany_bottom_in[100]}),
		.sram(mux_tree_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_59_sram_inv[0:1]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size2 mux_left_track_155 (
		.in({chany_top_in[37], chany_bottom_in[101]}),
		.sram(mux_tree_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_60_sram_inv[0:1]),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_size2 mux_left_track_157 (
		.in({chany_top_in[36], chany_bottom_in[102]}),
		.sram(mux_tree_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_61_sram_inv[0:1]),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_size2 mux_left_track_159 (
		.in({chany_top_in[34], chany_top_in[104]}),
		.sram(mux_tree_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_62_sram_inv[0:1]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_size2 mux_left_track_161 (
		.in({chany_top_in[33], chany_top_in[103]}),
		.sram(mux_tree_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_63_sram_inv[0:1]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size2 mux_left_track_165 (
		.in({chany_top_in[30], chany_top_in[95]}),
		.sram(mux_tree_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_64_sram_inv[0:1]),
		.out(chanx_left_out[82]));

	mux_tree_tapbuf_size2 mux_left_track_167 (
		.in({chany_top_in[29], chany_top_in[91]}),
		.sram(mux_tree_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_65_sram_inv[0:1]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_size2 mux_left_track_169 (
		.in({chany_top_in[28], chany_top_in[87]}),
		.sram(mux_tree_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_66_sram_inv[0:1]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size2 mux_left_track_171 (
		.in({chany_top_in[26], chany_top_in[83]}),
		.sram(mux_tree_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_67_sram_inv[0:1]),
		.out(chanx_left_out[85]));

	mux_tree_tapbuf_size2 mux_left_track_173 (
		.in({chany_top_in[25], chany_top_in[79]}),
		.sram(mux_tree_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_68_sram_inv[0:1]),
		.out(chanx_left_out[86]));

	mux_tree_tapbuf_size2 mux_left_track_175 (
		.in({chany_top_in[24], chany_top_in[75]}),
		.sram(mux_tree_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_69_sram_inv[0:1]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_size2 mux_left_track_177 (
		.in({chany_top_in[22], chany_top_in[71]}),
		.sram(mux_tree_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_70_sram_inv[0:1]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size2 mux_left_track_179 (
		.in({chany_top_in[21], chany_top_in[67]}),
		.sram(mux_tree_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_71_sram_inv[0:1]),
		.out(chanx_left_out[89]));

	mux_tree_tapbuf_size2 mux_left_track_185 (
		.in({chany_top_in[17], chany_top_in[55]}),
		.sram(mux_tree_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_72_sram_inv[0:1]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size2 mux_left_track_187 (
		.in({chany_top_in[16], chany_top_in[51]}),
		.sram(mux_tree_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_73_sram_inv[0:1]),
		.out(chanx_left_out[93]));

	mux_tree_tapbuf_size2 mux_left_track_189 (
		.in({chany_top_in[14], chany_top_in[47]}),
		.sram(mux_tree_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_74_sram_inv[0:1]),
		.out(chanx_left_out[94]));

	mux_tree_tapbuf_size2 mux_left_track_191 (
		.in({chany_top_in[13], chany_top_in[43]}),
		.sram(mux_tree_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_75_sram_inv[0:1]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_size2 mux_left_track_193 (
		.in({chany_top_in[12], chany_top_in[39]}),
		.sram(mux_tree_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_76_sram_inv[0:1]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size2 mux_left_track_195 (
		.in({chany_top_in[10], chany_top_in[35]}),
		.sram(mux_tree_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_77_sram_inv[0:1]),
		.out(chanx_left_out[97]));

	mux_tree_tapbuf_size2 mux_left_track_197 (
		.in({chany_top_in[9], chany_top_in[31]}),
		.sram(mux_tree_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_78_sram_inv[0:1]),
		.out(chanx_left_out[98]));

	mux_tree_tapbuf_size2 mux_left_track_201 (
		.in({chany_top_in[6], chany_top_in[23]}),
		.sram(mux_tree_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_79_sram_inv[0:1]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size2 mux_left_track_205 (
		.in({chany_top_in[4], chany_top_in[15]}),
		.sram(mux_tree_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_80_sram_inv[0:1]),
		.out(chanx_left_out[102]));

	mux_tree_tapbuf_size2 mux_left_track_207 (
		.in({chany_top_in[2], chany_top_in[11]}),
		.sram(mux_tree_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_81_sram_inv[0:1]),
		.out(chanx_left_out[103]));

	mux_tree_tapbuf_size2 mux_left_track_209 (
		.in({chany_top_in[1], chany_top_in[7]}),
		.sram(mux_tree_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_82_sram_inv[0:1]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size2_mem mem_left_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_27_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_28_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_29_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_30_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_31_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_32_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_33_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_34_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_35_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_36_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_37_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_38_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_39_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_40_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_41_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_42_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_43_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_44_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_45_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_46_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_47_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_48_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_49_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_50_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_51_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_52_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_53_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_54_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_55_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_147 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_56_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_149 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_57_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_151 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_58_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_59_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_155 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_60_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_157 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_61_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_159 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_62_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_63_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_165 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_64_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_167 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_65_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_66_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_171 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_67_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_173 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_68_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_175 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_69_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_70_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_179 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_71_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_72_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_187 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_73_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_189 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_74_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_191 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_75_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_76_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_195 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_77_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_197 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_78_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_79_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_205 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_80_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_207 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_81_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_82_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_10__3_ -----

//----- Default net type -----
`default_nettype wire



