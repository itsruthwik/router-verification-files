//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[4][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sat Jun 29 10:24:45 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_4__2_ -----
module sb_4__2_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_,
                ccff_head,
                chany_top_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:72] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:72] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
//----- INPUT PORTS -----
input [0:72] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:72] chany_top_out;
//----- OUTPUT PORTS -----
output [0:72] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:72] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size10_0_sram;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_1_sram;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail;
wire [0:3] mux_tree_tapbuf_size11_0_sram;
wire [0:3] mux_tree_tapbuf_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_10_sram;
wire [0:3] mux_tree_tapbuf_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_11_sram;
wire [0:3] mux_tree_tapbuf_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_12_sram;
wire [0:3] mux_tree_tapbuf_size11_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_1_sram;
wire [0:3] mux_tree_tapbuf_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_2_sram;
wire [0:3] mux_tree_tapbuf_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_3_sram;
wire [0:3] mux_tree_tapbuf_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_4_sram;
wire [0:3] mux_tree_tapbuf_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_5_sram;
wire [0:3] mux_tree_tapbuf_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_6_sram;
wire [0:3] mux_tree_tapbuf_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_7_sram;
wire [0:3] mux_tree_tapbuf_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_8_sram;
wire [0:3] mux_tree_tapbuf_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_9_sram;
wire [0:3] mux_tree_tapbuf_size11_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size12_0_sram;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_10_sram;
wire [0:3] mux_tree_tapbuf_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_11_sram;
wire [0:3] mux_tree_tapbuf_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_12_sram;
wire [0:3] mux_tree_tapbuf_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_13_sram;
wire [0:3] mux_tree_tapbuf_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_14_sram;
wire [0:3] mux_tree_tapbuf_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_15_sram;
wire [0:3] mux_tree_tapbuf_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_16_sram;
wire [0:3] mux_tree_tapbuf_size12_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_17_sram;
wire [0:3] mux_tree_tapbuf_size12_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_18_sram;
wire [0:3] mux_tree_tapbuf_size12_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_19_sram;
wire [0:3] mux_tree_tapbuf_size12_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_1_sram;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_20_sram;
wire [0:3] mux_tree_tapbuf_size12_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_21_sram;
wire [0:3] mux_tree_tapbuf_size12_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_22_sram;
wire [0:3] mux_tree_tapbuf_size12_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_23_sram;
wire [0:3] mux_tree_tapbuf_size12_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_24_sram;
wire [0:3] mux_tree_tapbuf_size12_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_25_sram;
wire [0:3] mux_tree_tapbuf_size12_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_26_sram;
wire [0:3] mux_tree_tapbuf_size12_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_27_sram;
wire [0:3] mux_tree_tapbuf_size12_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_28_sram;
wire [0:3] mux_tree_tapbuf_size12_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_29_sram;
wire [0:3] mux_tree_tapbuf_size12_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_2_sram;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_30_sram;
wire [0:3] mux_tree_tapbuf_size12_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_31_sram;
wire [0:3] mux_tree_tapbuf_size12_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_32_sram;
wire [0:3] mux_tree_tapbuf_size12_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_33_sram;
wire [0:3] mux_tree_tapbuf_size12_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_34_sram;
wire [0:3] mux_tree_tapbuf_size12_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_35_sram;
wire [0:3] mux_tree_tapbuf_size12_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_36_sram;
wire [0:3] mux_tree_tapbuf_size12_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_37_sram;
wire [0:3] mux_tree_tapbuf_size12_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_38_sram;
wire [0:3] mux_tree_tapbuf_size12_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_39_sram;
wire [0:3] mux_tree_tapbuf_size12_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_3_sram;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_40_sram;
wire [0:3] mux_tree_tapbuf_size12_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_4_sram;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_5_sram;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_6_sram;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_7_sram;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_8_sram;
wire [0:3] mux_tree_tapbuf_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_9_sram;
wire [0:3] mux_tree_tapbuf_size12_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size13_0_sram;
wire [0:3] mux_tree_tapbuf_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_10_sram;
wire [0:3] mux_tree_tapbuf_size13_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_11_sram;
wire [0:3] mux_tree_tapbuf_size13_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_12_sram;
wire [0:3] mux_tree_tapbuf_size13_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_13_sram;
wire [0:3] mux_tree_tapbuf_size13_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_14_sram;
wire [0:3] mux_tree_tapbuf_size13_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_15_sram;
wire [0:3] mux_tree_tapbuf_size13_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_1_sram;
wire [0:3] mux_tree_tapbuf_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_2_sram;
wire [0:3] mux_tree_tapbuf_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_3_sram;
wire [0:3] mux_tree_tapbuf_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_4_sram;
wire [0:3] mux_tree_tapbuf_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_5_sram;
wire [0:3] mux_tree_tapbuf_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_6_sram;
wire [0:3] mux_tree_tapbuf_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_7_sram;
wire [0:3] mux_tree_tapbuf_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_8_sram;
wire [0:3] mux_tree_tapbuf_size13_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_9_sram;
wire [0:3] mux_tree_tapbuf_size13_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size14_0_sram;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail;
wire [0:4] mux_tree_tapbuf_size20_0_sram;
wire [0:4] mux_tree_tapbuf_size20_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_1_sram;
wire [0:4] mux_tree_tapbuf_size20_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_2_sram;
wire [0:4] mux_tree_tapbuf_size20_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_3_sram;
wire [0:4] mux_tree_tapbuf_size20_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_4_sram;
wire [0:4] mux_tree_tapbuf_size20_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_5_sram;
wire [0:4] mux_tree_tapbuf_size20_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_6_sram;
wire [0:4] mux_tree_tapbuf_size20_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_7_sram;
wire [0:4] mux_tree_tapbuf_size20_7_sram_inv;
wire [0:0] mux_tree_tapbuf_size20_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_7_ccff_tail;
wire [0:4] mux_tree_tapbuf_size21_0_sram;
wire [0:4] mux_tree_tapbuf_size21_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_1_sram;
wire [0:4] mux_tree_tapbuf_size21_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_2_sram;
wire [0:4] mux_tree_tapbuf_size21_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_3_sram;
wire [0:4] mux_tree_tapbuf_size21_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_4_sram;
wire [0:4] mux_tree_tapbuf_size21_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_5_sram;
wire [0:4] mux_tree_tapbuf_size21_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_6_sram;
wire [0:4] mux_tree_tapbuf_size21_6_sram_inv;
wire [0:0] mux_tree_tapbuf_size21_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_6_ccff_tail;
wire [0:4] mux_tree_tapbuf_size22_0_sram;
wire [0:4] mux_tree_tapbuf_size22_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size22_1_sram;
wire [0:4] mux_tree_tapbuf_size22_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size22_2_sram;
wire [0:4] mux_tree_tapbuf_size22_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size22_3_sram;
wire [0:4] mux_tree_tapbuf_size22_3_sram_inv;
wire [0:0] mux_tree_tapbuf_size22_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size22_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size22_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size22_mem_3_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size7 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[0], chanx_left_in[19], chanx_left_in[38], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size7 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[12], chanx_left_in[31], chanx_left_in[50], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size7_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[18], chanx_left_in[37], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size6 mux_top_track_32 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[15], chanx_left_in[34], chanx_left_in[53], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size6 mux_top_track_40 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[14], chanx_left_in[33], chanx_left_in[52], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size6 mux_top_track_48 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[13], chanx_left_in[32], chanx_left_in[51], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size6 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[11], chanx_left_in[30], chanx_left_in[49], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size6 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[10], chanx_left_in[29], chanx_left_in[48], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size6 mux_top_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[6], chanx_left_in[25], chanx_left_in[44], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size6 mux_top_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[5], chanx_left_in[24], chanx_left_in[43], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size6 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[1], chanx_left_in[20], chanx_left_in[39], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size6_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[17], chanx_left_in[36], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size5 mux_top_track_24 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[16], chanx_left_in[35], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size5 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[9], chanx_left_in[28], chanx_left_in[47], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size5 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[8], chanx_left_in[27], chanx_left_in[46], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size5 mux_top_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[7], chanx_left_in[26], chanx_left_in[45], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size5 mux_top_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[4], chanx_left_in[23], chanx_left_in[42], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size5 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[3], chanx_left_in[22], chanx_left_in[41], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size5 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[2], chanx_left_in[21], chanx_left_in[40], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size5_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size22 mux_bottom_track_1 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[1], chanx_left_in[20], chanx_left_in[39], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_size22_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_0_sram_inv[0:4]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size22 mux_bottom_track_49 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[7], chanx_left_in[26], chanx_left_in[45], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_size22_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_1_sram_inv[0:4]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size22 mux_bottom_track_57 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[8], chanx_left_in[27], chanx_left_in[46], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_size22_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_2_sram_inv[0:4]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size22 mux_bottom_track_145 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[0], chanx_left_in[19], chanx_left_in[38], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_size22_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_3_sram_inv[0:4]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size22_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_0_sram_inv[0:4]));

	mux_tree_tapbuf_size22_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_1_sram_inv[0:4]));

	mux_tree_tapbuf_size22_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_2_sram_inv[0:4]));

	mux_tree_tapbuf_size22_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_3_sram_inv[0:4]));

	mux_tree_tapbuf_size21 mux_bottom_track_9 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[2], chanx_left_in[21], chanx_left_in[40], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_size21_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_0_sram_inv[0:4]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size21 mux_bottom_track_41 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[6], chanx_left_in[25], chanx_left_in[44], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_size21_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_1_sram_inv[0:4]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size21 mux_bottom_track_65 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[9], chanx_left_in[28], chanx_left_in[47], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_size21_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_2_sram_inv[0:4]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size21 mux_bottom_track_73 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[10], chanx_left_in[29], chanx_left_in[48], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_size21_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_3_sram_inv[0:4]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size21 mux_bottom_track_97 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[13], chanx_left_in[32], chanx_left_in[51], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_size21_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_4_sram_inv[0:4]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size21 mux_bottom_track_105 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[14], chanx_left_in[33], chanx_left_in[52], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_size21_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_5_sram_inv[0:4]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size21 mux_bottom_track_113 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[15], chanx_left_in[34], chanx_left_in[53], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_size21_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_6_sram_inv[0:4]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_0_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_1_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_2_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_3_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_4_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_5_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_6_sram_inv[0:4]));

	mux_tree_tapbuf_size20 mux_bottom_track_17 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[3], chanx_left_in[22], chanx_left_in[41], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_size20_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_0_sram_inv[0:4]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size20 mux_bottom_track_25 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[4], chanx_left_in[23], chanx_left_in[42], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_size20_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_1_sram_inv[0:4]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size20 mux_bottom_track_33 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[5], chanx_left_in[24], chanx_left_in[43], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_size20_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_2_sram_inv[0:4]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size20 mux_bottom_track_81 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[11], chanx_left_in[30], chanx_left_in[49], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_size20_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_3_sram_inv[0:4]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size20 mux_bottom_track_89 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[12], chanx_left_in[31], chanx_left_in[50], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_size20_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_4_sram_inv[0:4]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size20 mux_bottom_track_121 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[16], chanx_left_in[35], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_size20_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_5_sram_inv[0:4]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size20 mux_bottom_track_129 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[17], chanx_left_in[36], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_size20_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_6_sram_inv[0:4]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size20 mux_bottom_track_137 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[18], chanx_left_in[37], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_size20_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_7_sram_inv[0:4]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_0_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_1_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_2_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_3_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_4_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_5_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_6_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_7_sram_inv[0:4]));

	mux_tree_tapbuf_size12 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_0_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size12 mux_left_track_5 (
		.in({chany_bottom_in[1], chany_bottom_in[7], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_1_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_size12 mux_left_track_15 (
		.in({chany_bottom_in[8], chany_bottom_in[27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_2_sram_inv[0:3]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_size12 mux_left_track_17 (
		.in({chany_bottom_in[9], chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_3_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size12 mux_left_track_21 (
		.in({chany_bottom_in[12], chany_bottom_in[39], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_4_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_size12 mux_left_track_31 (
		.in({chany_bottom_in[18], chany_bottom_in[59], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_5_sram_inv[0:3]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_size12 mux_left_track_37 (
		.in({chany_bottom_in[22], chany_bottom_in[71], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_6_sram_inv[0:3]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_size12 mux_left_track_39 (
		.in({chany_bottom_in[24], chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_7_sram_inv[0:3]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_size12 mux_left_track_41 (
		.in({chany_top_in[70], chany_bottom_in[25], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_8_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size12 mux_left_track_43 (
		.in({chany_top_in[69], chany_bottom_in[26], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_9_sram_inv[0:3]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_size12 mux_left_track_47 (
		.in({chany_top_in[66], chany_bottom_in[29], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_10_sram_inv[0:3]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_size12 mux_left_track_55 (
		.in({chany_top_in[61], chany_bottom_in[34], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_11_sram_inv[0:3]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_size12 mux_left_track_57 (
		.in({chany_top_in[60], chany_bottom_in[36], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_12_sram_inv[0:3]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size12 mux_left_track_59 (
		.in({chany_top_in[58], chany_bottom_in[37], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_13_sram_inv[0:3]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_size12 mux_left_track_61 (
		.in({chany_top_in[57], chany_bottom_in[38], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_14_sram_inv[0:3]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_size12 mux_left_track_65 (
		.in({chany_top_in[54], chany_bottom_in[41], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_15_sram_inv[0:3]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size12 mux_left_track_69 (
		.in({chany_top_in[52], chany_bottom_in[44], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_16_sram_inv[0:3]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_size12 mux_left_track_73 (
		.in({chany_top_in[49], chany_bottom_in[46], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_17_sram_inv[0:3]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size12 mux_left_track_75 (
		.in({chany_top_in[48], chany_bottom_in[48], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_18_sram_inv[0:3]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_size12 mux_left_track_77 (
		.in({chany_top_in[46], chany_bottom_in[49], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_19_sram_inv[0:3]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_size12 mux_left_track_79 (
		.in({chany_top_in[45], chany_bottom_in[50], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_20_sram_inv[0:3]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_size12 mux_left_track_83 (
		.in({chany_top_in[42], chany_bottom_in[53], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_21_sram_inv[0:3]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_size12 mux_left_track_85 (
		.in({chany_top_in[41], chany_bottom_in[54], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_22_sram_inv[0:3]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_size12 mux_left_track_93 (
		.in({chany_top_in[36], chany_bottom_in[60], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_23_sram_inv[0:3]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_size12 mux_left_track_95 (
		.in({chany_top_in[34], chany_bottom_in[61], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_24_sram_inv[0:3]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_size12 mux_left_track_97 (
		.in({chany_top_in[33], chany_bottom_in[62], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_25_sram_inv[0:3]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size12 mux_left_track_101 (
		.in({chany_top_in[30], chany_bottom_in[65], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_26_sram_inv[0:3]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_size12 mux_left_track_103 (
		.in({chany_top_in[29], chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_27_sram_inv[0:3]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_size12 mux_left_track_105 (
		.in({chany_top_in[28], chany_bottom_in[68], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_28_sram_inv[0:3]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size12 mux_left_track_109 (
		.in({chany_top_in[25], chany_bottom_in[70], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_29_sram_inv[0:3]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_size12 mux_left_track_113 (
		.in({chany_top_in[22], chany_top_in[71], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_30_sram_inv[0:3]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size12 mux_left_track_115 (
		.in({chany_top_in[21], chany_top_in[67], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_31_sram_inv[0:3]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_size12 mux_left_track_119 (
		.in({chany_top_in[18], chany_top_in[59], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_32_sram_inv[0:3]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_size12 mux_left_track_121 (
		.in({chany_top_in[17], chany_top_in[55], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_33_sram_inv[0:3]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size12 mux_left_track_123 (
		.in({chany_top_in[16], chany_top_in[51], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_34_sram_inv[0:3]),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_size12 mux_left_track_129 (
		.in({chany_top_in[12], chany_top_in[39], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_35_sram_inv[0:3]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size12 mux_left_track_133 (
		.in({chany_top_in[9], chany_top_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_36_sram_inv[0:3]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_size12 mux_left_track_137 (
		.in({chany_top_in[6], chany_top_in[23], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_37_sram_inv[0:3]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size12 mux_left_track_139 (
		.in({chany_top_in[5], chany_top_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_38_sram_inv[0:3]),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_size12 mux_left_track_141 (
		.in({chany_top_in[4], chany_top_in[15], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_39_sram_inv[0:3]),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_size12 mux_left_track_145 (
		.in({chany_top_in[1], chany_top_in[7], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_40_sram_inv[0:3]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size12_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_16_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_17_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_18_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_19_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_20_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_21_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_22_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_23_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_24_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_25_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_26_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_27_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_28_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_29_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_30_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_31_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_32_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_33_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_34_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_35_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_36_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_37_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_38_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_39_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_40_sram_inv[0:3]));

	mux_tree_tapbuf_size13 mux_left_track_3 (
		.in({chany_bottom_in[0], chany_bottom_in[3], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_0_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_size13 mux_left_track_9 (
		.in({chany_bottom_in[4], chany_bottom_in[15], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_1_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size13 mux_left_track_11 (
		.in({chany_bottom_in[5], chany_bottom_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_2_sram_inv[0:3]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_size13 mux_left_track_13 (
		.in({chany_bottom_in[6], chany_bottom_in[23], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_3_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_size13 mux_left_track_19 (
		.in({chany_bottom_in[10], chany_bottom_in[35], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_4_sram_inv[0:3]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_size13 mux_left_track_23 (
		.in({chany_bottom_in[13], chany_bottom_in[43], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_5_sram_inv[0:3]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_size13 mux_left_track_25 (
		.in({chany_bottom_in[14], chany_bottom_in[47], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_6_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size13 mux_left_track_27 (
		.in({chany_bottom_in[16], chany_bottom_in[51], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_7_sram_inv[0:3]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_size13 mux_left_track_29 (
		.in({chany_bottom_in[17], chany_bottom_in[55], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_8_sram_inv[0:3]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_size13 mux_left_track_45 (
		.in({chany_top_in[68], chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_9_sram_inv[0:3]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_size13 mux_left_track_49 (
		.in({chany_top_in[65], chany_bottom_in[30], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size13_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_10_sram_inv[0:3]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size13 mux_left_track_63 (
		.in({chany_top_in[56], chany_bottom_in[40], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_11_sram_inv[0:3]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_size13 mux_left_track_81 (
		.in({chany_top_in[44], chany_bottom_in[52], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_12_sram_inv[0:3]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size13 mux_left_track_99 (
		.in({chany_top_in[32], chany_bottom_in[64], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_13_sram_inv[0:3]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_size13 mux_left_track_117 (
		.in({chany_top_in[20], chany_top_in[63], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_14_sram_inv[0:3]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_size13 mux_left_track_135 (
		.in({chany_top_in[8], chany_top_in[27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_15_sram_inv[0:3]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_size13_mem mem_left_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_9_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_10_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_11_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_12_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_13_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_14_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_15_sram_inv[0:3]));

	mux_tree_tapbuf_size14 mux_left_track_7 (
		.in({chany_bottom_in[2], chany_bottom_in[11], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size14_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_0_sram_inv[0:3]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_size14_mem mem_left_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11 mux_left_track_33 (
		.in({chany_bottom_in[20], chany_bottom_in[63], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_0_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size11 mux_left_track_35 (
		.in({chany_bottom_in[21], chany_bottom_in[67], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_1_sram_inv[0:3]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_size11 mux_left_track_51 (
		.in({chany_top_in[64], chany_bottom_in[32], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_2_sram_inv[0:3]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_size11 mux_left_track_53 (
		.in({chany_top_in[62], chany_bottom_in[33], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_3_sram_inv[0:3]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_size11 mux_left_track_67 (
		.in({chany_top_in[53], chany_bottom_in[42], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_4_sram_inv[0:3]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_size11 mux_left_track_87 (
		.in({chany_top_in[40], chany_bottom_in[56], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_5_sram_inv[0:3]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_size11 mux_left_track_89 (
		.in({chany_top_in[38], chany_bottom_in[57], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_6_sram_inv[0:3]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size11 mux_left_track_91 (
		.in({chany_top_in[37], chany_bottom_in[58], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_7_sram_inv[0:3]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_size11 mux_left_track_111 (
		.in({chany_top_in[24], chany_top_in[72], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_8_sram_inv[0:3]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_size11 mux_left_track_125 (
		.in({chany_top_in[14], chany_top_in[47], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_9_sram_inv[0:3]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_size11 mux_left_track_127 (
		.in({chany_top_in[13], chany_top_in[43], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_10_sram_inv[0:3]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_size11 mux_left_track_131 (
		.in({chany_top_in[10], chany_top_in[35], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_11_sram_inv[0:3]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_size11 mux_left_track_143 (
		.in({chany_top_in[2], chany_top_in[11], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size11_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_12_sram_inv[0:3]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_size11_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_12_sram_inv[0:3]));

	mux_tree_tapbuf_size10 mux_left_track_71 (
		.in({chany_top_in[50], chany_bottom_in[45], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_0_sram_inv[0:3]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_size10 mux_left_track_107 (
		.in({chany_top_in[26], chany_bottom_in[69], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_1_sram_inv[0:3]),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_size10_mem mem_left_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_1_sram_inv[0:3]));

endmodule
// ----- END Verilog module for sb_4__2_ -----

//----- Default net type -----
`default_nettype wire



