//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[4][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jun 28 12:51:27 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_4__1_ -----
module sb_4__1_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                ccff_head,
                chany_top_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:192] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:192] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:192] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:192] chany_top_out;
//----- OUTPUT PORTS -----
output [0:192] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:192] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size10_0_sram;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_10_sram;
wire [0:3] mux_tree_tapbuf_size10_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_11_sram;
wire [0:3] mux_tree_tapbuf_size10_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_12_sram;
wire [0:3] mux_tree_tapbuf_size10_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_13_sram;
wire [0:3] mux_tree_tapbuf_size10_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_14_sram;
wire [0:3] mux_tree_tapbuf_size10_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_15_sram;
wire [0:3] mux_tree_tapbuf_size10_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_16_sram;
wire [0:3] mux_tree_tapbuf_size10_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_1_sram;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_2_sram;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_3_sram;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_4_sram;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_5_sram;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_6_sram;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_7_sram;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_8_sram;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_9_sram;
wire [0:3] mux_tree_tapbuf_size10_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size11_0_sram;
wire [0:3] mux_tree_tapbuf_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_10_sram;
wire [0:3] mux_tree_tapbuf_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_11_sram;
wire [0:3] mux_tree_tapbuf_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_12_sram;
wire [0:3] mux_tree_tapbuf_size11_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_13_sram;
wire [0:3] mux_tree_tapbuf_size11_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_14_sram;
wire [0:3] mux_tree_tapbuf_size11_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_15_sram;
wire [0:3] mux_tree_tapbuf_size11_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_16_sram;
wire [0:3] mux_tree_tapbuf_size11_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_17_sram;
wire [0:3] mux_tree_tapbuf_size11_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_18_sram;
wire [0:3] mux_tree_tapbuf_size11_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_19_sram;
wire [0:3] mux_tree_tapbuf_size11_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_1_sram;
wire [0:3] mux_tree_tapbuf_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_20_sram;
wire [0:3] mux_tree_tapbuf_size11_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_21_sram;
wire [0:3] mux_tree_tapbuf_size11_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_22_sram;
wire [0:3] mux_tree_tapbuf_size11_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_23_sram;
wire [0:3] mux_tree_tapbuf_size11_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_24_sram;
wire [0:3] mux_tree_tapbuf_size11_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_25_sram;
wire [0:3] mux_tree_tapbuf_size11_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_26_sram;
wire [0:3] mux_tree_tapbuf_size11_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_27_sram;
wire [0:3] mux_tree_tapbuf_size11_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_28_sram;
wire [0:3] mux_tree_tapbuf_size11_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_29_sram;
wire [0:3] mux_tree_tapbuf_size11_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_2_sram;
wire [0:3] mux_tree_tapbuf_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_30_sram;
wire [0:3] mux_tree_tapbuf_size11_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_31_sram;
wire [0:3] mux_tree_tapbuf_size11_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_32_sram;
wire [0:3] mux_tree_tapbuf_size11_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_33_sram;
wire [0:3] mux_tree_tapbuf_size11_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_34_sram;
wire [0:3] mux_tree_tapbuf_size11_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_35_sram;
wire [0:3] mux_tree_tapbuf_size11_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_36_sram;
wire [0:3] mux_tree_tapbuf_size11_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_37_sram;
wire [0:3] mux_tree_tapbuf_size11_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_38_sram;
wire [0:3] mux_tree_tapbuf_size11_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_39_sram;
wire [0:3] mux_tree_tapbuf_size11_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_3_sram;
wire [0:3] mux_tree_tapbuf_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_40_sram;
wire [0:3] mux_tree_tapbuf_size11_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_41_sram;
wire [0:3] mux_tree_tapbuf_size11_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_42_sram;
wire [0:3] mux_tree_tapbuf_size11_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_43_sram;
wire [0:3] mux_tree_tapbuf_size11_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_44_sram;
wire [0:3] mux_tree_tapbuf_size11_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_45_sram;
wire [0:3] mux_tree_tapbuf_size11_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_46_sram;
wire [0:3] mux_tree_tapbuf_size11_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_47_sram;
wire [0:3] mux_tree_tapbuf_size11_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_48_sram;
wire [0:3] mux_tree_tapbuf_size11_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_49_sram;
wire [0:3] mux_tree_tapbuf_size11_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_4_sram;
wire [0:3] mux_tree_tapbuf_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_50_sram;
wire [0:3] mux_tree_tapbuf_size11_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_51_sram;
wire [0:3] mux_tree_tapbuf_size11_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_52_sram;
wire [0:3] mux_tree_tapbuf_size11_52_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_53_sram;
wire [0:3] mux_tree_tapbuf_size11_53_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_54_sram;
wire [0:3] mux_tree_tapbuf_size11_54_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_55_sram;
wire [0:3] mux_tree_tapbuf_size11_55_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_56_sram;
wire [0:3] mux_tree_tapbuf_size11_56_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_57_sram;
wire [0:3] mux_tree_tapbuf_size11_57_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_58_sram;
wire [0:3] mux_tree_tapbuf_size11_58_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_59_sram;
wire [0:3] mux_tree_tapbuf_size11_59_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_5_sram;
wire [0:3] mux_tree_tapbuf_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_60_sram;
wire [0:3] mux_tree_tapbuf_size11_60_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_61_sram;
wire [0:3] mux_tree_tapbuf_size11_61_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_62_sram;
wire [0:3] mux_tree_tapbuf_size11_62_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_63_sram;
wire [0:3] mux_tree_tapbuf_size11_63_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_64_sram;
wire [0:3] mux_tree_tapbuf_size11_64_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_65_sram;
wire [0:3] mux_tree_tapbuf_size11_65_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_66_sram;
wire [0:3] mux_tree_tapbuf_size11_66_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_67_sram;
wire [0:3] mux_tree_tapbuf_size11_67_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_68_sram;
wire [0:3] mux_tree_tapbuf_size11_68_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_69_sram;
wire [0:3] mux_tree_tapbuf_size11_69_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_6_sram;
wire [0:3] mux_tree_tapbuf_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_70_sram;
wire [0:3] mux_tree_tapbuf_size11_70_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_71_sram;
wire [0:3] mux_tree_tapbuf_size11_71_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_7_sram;
wire [0:3] mux_tree_tapbuf_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_8_sram;
wire [0:3] mux_tree_tapbuf_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_9_sram;
wire [0:3] mux_tree_tapbuf_size11_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size12_0_sram;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_10_sram;
wire [0:3] mux_tree_tapbuf_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_11_sram;
wire [0:3] mux_tree_tapbuf_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_12_sram;
wire [0:3] mux_tree_tapbuf_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_13_sram;
wire [0:3] mux_tree_tapbuf_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_14_sram;
wire [0:3] mux_tree_tapbuf_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_15_sram;
wire [0:3] mux_tree_tapbuf_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_16_sram;
wire [0:3] mux_tree_tapbuf_size12_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_17_sram;
wire [0:3] mux_tree_tapbuf_size12_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_18_sram;
wire [0:3] mux_tree_tapbuf_size12_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_19_sram;
wire [0:3] mux_tree_tapbuf_size12_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_1_sram;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_20_sram;
wire [0:3] mux_tree_tapbuf_size12_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_21_sram;
wire [0:3] mux_tree_tapbuf_size12_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_22_sram;
wire [0:3] mux_tree_tapbuf_size12_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_23_sram;
wire [0:3] mux_tree_tapbuf_size12_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_24_sram;
wire [0:3] mux_tree_tapbuf_size12_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_25_sram;
wire [0:3] mux_tree_tapbuf_size12_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_26_sram;
wire [0:3] mux_tree_tapbuf_size12_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_27_sram;
wire [0:3] mux_tree_tapbuf_size12_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_28_sram;
wire [0:3] mux_tree_tapbuf_size12_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_29_sram;
wire [0:3] mux_tree_tapbuf_size12_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_2_sram;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_30_sram;
wire [0:3] mux_tree_tapbuf_size12_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_31_sram;
wire [0:3] mux_tree_tapbuf_size12_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_32_sram;
wire [0:3] mux_tree_tapbuf_size12_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_33_sram;
wire [0:3] mux_tree_tapbuf_size12_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_34_sram;
wire [0:3] mux_tree_tapbuf_size12_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_35_sram;
wire [0:3] mux_tree_tapbuf_size12_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_36_sram;
wire [0:3] mux_tree_tapbuf_size12_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_37_sram;
wire [0:3] mux_tree_tapbuf_size12_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_38_sram;
wire [0:3] mux_tree_tapbuf_size12_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_39_sram;
wire [0:3] mux_tree_tapbuf_size12_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_3_sram;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_40_sram;
wire [0:3] mux_tree_tapbuf_size12_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_41_sram;
wire [0:3] mux_tree_tapbuf_size12_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_42_sram;
wire [0:3] mux_tree_tapbuf_size12_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_43_sram;
wire [0:3] mux_tree_tapbuf_size12_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_44_sram;
wire [0:3] mux_tree_tapbuf_size12_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_45_sram;
wire [0:3] mux_tree_tapbuf_size12_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_46_sram;
wire [0:3] mux_tree_tapbuf_size12_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_47_sram;
wire [0:3] mux_tree_tapbuf_size12_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_48_sram;
wire [0:3] mux_tree_tapbuf_size12_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_49_sram;
wire [0:3] mux_tree_tapbuf_size12_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_4_sram;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_50_sram;
wire [0:3] mux_tree_tapbuf_size12_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_51_sram;
wire [0:3] mux_tree_tapbuf_size12_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_52_sram;
wire [0:3] mux_tree_tapbuf_size12_52_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_53_sram;
wire [0:3] mux_tree_tapbuf_size12_53_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_54_sram;
wire [0:3] mux_tree_tapbuf_size12_54_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_55_sram;
wire [0:3] mux_tree_tapbuf_size12_55_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_56_sram;
wire [0:3] mux_tree_tapbuf_size12_56_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_57_sram;
wire [0:3] mux_tree_tapbuf_size12_57_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_58_sram;
wire [0:3] mux_tree_tapbuf_size12_58_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_59_sram;
wire [0:3] mux_tree_tapbuf_size12_59_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_5_sram;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_60_sram;
wire [0:3] mux_tree_tapbuf_size12_60_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_61_sram;
wire [0:3] mux_tree_tapbuf_size12_61_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_62_sram;
wire [0:3] mux_tree_tapbuf_size12_62_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_63_sram;
wire [0:3] mux_tree_tapbuf_size12_63_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_64_sram;
wire [0:3] mux_tree_tapbuf_size12_64_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_65_sram;
wire [0:3] mux_tree_tapbuf_size12_65_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_66_sram;
wire [0:3] mux_tree_tapbuf_size12_66_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_67_sram;
wire [0:3] mux_tree_tapbuf_size12_67_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_68_sram;
wire [0:3] mux_tree_tapbuf_size12_68_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_69_sram;
wire [0:3] mux_tree_tapbuf_size12_69_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_6_sram;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_70_sram;
wire [0:3] mux_tree_tapbuf_size12_70_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_71_sram;
wire [0:3] mux_tree_tapbuf_size12_71_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_72_sram;
wire [0:3] mux_tree_tapbuf_size12_72_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_73_sram;
wire [0:3] mux_tree_tapbuf_size12_73_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_74_sram;
wire [0:3] mux_tree_tapbuf_size12_74_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_75_sram;
wire [0:3] mux_tree_tapbuf_size12_75_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_76_sram;
wire [0:3] mux_tree_tapbuf_size12_76_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_77_sram;
wire [0:3] mux_tree_tapbuf_size12_77_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_78_sram;
wire [0:3] mux_tree_tapbuf_size12_78_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_79_sram;
wire [0:3] mux_tree_tapbuf_size12_79_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_7_sram;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_80_sram;
wire [0:3] mux_tree_tapbuf_size12_80_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_81_sram;
wire [0:3] mux_tree_tapbuf_size12_81_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_82_sram;
wire [0:3] mux_tree_tapbuf_size12_82_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_83_sram;
wire [0:3] mux_tree_tapbuf_size12_83_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_84_sram;
wire [0:3] mux_tree_tapbuf_size12_84_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_85_sram;
wire [0:3] mux_tree_tapbuf_size12_85_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_86_sram;
wire [0:3] mux_tree_tapbuf_size12_86_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_87_sram;
wire [0:3] mux_tree_tapbuf_size12_87_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_88_sram;
wire [0:3] mux_tree_tapbuf_size12_88_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_89_sram;
wire [0:3] mux_tree_tapbuf_size12_89_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_8_sram;
wire [0:3] mux_tree_tapbuf_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_9_sram;
wire [0:3] mux_tree_tapbuf_size12_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size13_0_sram;
wire [0:3] mux_tree_tapbuf_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_10_sram;
wire [0:3] mux_tree_tapbuf_size13_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_11_sram;
wire [0:3] mux_tree_tapbuf_size13_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_12_sram;
wire [0:3] mux_tree_tapbuf_size13_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_1_sram;
wire [0:3] mux_tree_tapbuf_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_2_sram;
wire [0:3] mux_tree_tapbuf_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_3_sram;
wire [0:3] mux_tree_tapbuf_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_4_sram;
wire [0:3] mux_tree_tapbuf_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_5_sram;
wire [0:3] mux_tree_tapbuf_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_6_sram;
wire [0:3] mux_tree_tapbuf_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_7_sram;
wire [0:3] mux_tree_tapbuf_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_8_sram;
wire [0:3] mux_tree_tapbuf_size13_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_9_sram;
wire [0:3] mux_tree_tapbuf_size13_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size15_0_sram;
wire [0:3] mux_tree_tapbuf_size15_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_1_sram;
wire [0:3] mux_tree_tapbuf_size15_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_2_sram;
wire [0:3] mux_tree_tapbuf_size15_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size15_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_2_ccff_tail;
wire [0:4] mux_tree_tapbuf_size16_0_sram;
wire [0:4] mux_tree_tapbuf_size16_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_10_sram;
wire [0:4] mux_tree_tapbuf_size16_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_11_sram;
wire [0:4] mux_tree_tapbuf_size16_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_12_sram;
wire [0:4] mux_tree_tapbuf_size16_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_13_sram;
wire [0:4] mux_tree_tapbuf_size16_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_14_sram;
wire [0:4] mux_tree_tapbuf_size16_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_15_sram;
wire [0:4] mux_tree_tapbuf_size16_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_16_sram;
wire [0:4] mux_tree_tapbuf_size16_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_17_sram;
wire [0:4] mux_tree_tapbuf_size16_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_18_sram;
wire [0:4] mux_tree_tapbuf_size16_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_19_sram;
wire [0:4] mux_tree_tapbuf_size16_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_1_sram;
wire [0:4] mux_tree_tapbuf_size16_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_20_sram;
wire [0:4] mux_tree_tapbuf_size16_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_21_sram;
wire [0:4] mux_tree_tapbuf_size16_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_22_sram;
wire [0:4] mux_tree_tapbuf_size16_22_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_23_sram;
wire [0:4] mux_tree_tapbuf_size16_23_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_24_sram;
wire [0:4] mux_tree_tapbuf_size16_24_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_25_sram;
wire [0:4] mux_tree_tapbuf_size16_25_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_2_sram;
wire [0:4] mux_tree_tapbuf_size16_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_3_sram;
wire [0:4] mux_tree_tapbuf_size16_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_4_sram;
wire [0:4] mux_tree_tapbuf_size16_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_5_sram;
wire [0:4] mux_tree_tapbuf_size16_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_6_sram;
wire [0:4] mux_tree_tapbuf_size16_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_7_sram;
wire [0:4] mux_tree_tapbuf_size16_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_8_sram;
wire [0:4] mux_tree_tapbuf_size16_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_9_sram;
wire [0:4] mux_tree_tapbuf_size16_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size16_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size17_0_sram;
wire [0:4] mux_tree_tapbuf_size17_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_10_sram;
wire [0:4] mux_tree_tapbuf_size17_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_11_sram;
wire [0:4] mux_tree_tapbuf_size17_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_12_sram;
wire [0:4] mux_tree_tapbuf_size17_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_13_sram;
wire [0:4] mux_tree_tapbuf_size17_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_14_sram;
wire [0:4] mux_tree_tapbuf_size17_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_15_sram;
wire [0:4] mux_tree_tapbuf_size17_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_16_sram;
wire [0:4] mux_tree_tapbuf_size17_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_17_sram;
wire [0:4] mux_tree_tapbuf_size17_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_1_sram;
wire [0:4] mux_tree_tapbuf_size17_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_2_sram;
wire [0:4] mux_tree_tapbuf_size17_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_3_sram;
wire [0:4] mux_tree_tapbuf_size17_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_4_sram;
wire [0:4] mux_tree_tapbuf_size17_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_5_sram;
wire [0:4] mux_tree_tapbuf_size17_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_6_sram;
wire [0:4] mux_tree_tapbuf_size17_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_7_sram;
wire [0:4] mux_tree_tapbuf_size17_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_8_sram;
wire [0:4] mux_tree_tapbuf_size17_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_9_sram;
wire [0:4] mux_tree_tapbuf_size17_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size17_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size18_0_sram;
wire [0:4] mux_tree_tapbuf_size18_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_1_sram;
wire [0:4] mux_tree_tapbuf_size18_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size18_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_1_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_29_sram;
wire [0:2] mux_tree_tapbuf_size5_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_30_sram;
wire [0:2] mux_tree_tapbuf_size5_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_31_sram;
wire [0:2] mux_tree_tapbuf_size5_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_32_sram;
wire [0:2] mux_tree_tapbuf_size5_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_33_sram;
wire [0:2] mux_tree_tapbuf_size5_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_10_sram;
wire [0:2] mux_tree_tapbuf_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_9_sram;
wire [0:2] mux_tree_tapbuf_size6_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:3] mux_tree_tapbuf_size9_0_sram;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[189] = chany_top_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[190] = chany_top_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[191] = chany_top_in[190];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[189] = chany_bottom_in[188];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[190] = chany_bottom_in[189];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[191] = chany_bottom_in[190];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size17 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[0], chanx_left_in[49], chanx_left_in[98], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size17_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_0_sram_inv[0:4]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size17 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[45], chanx_left_in[94], chanx_left_in[143], chanx_left_in[192]}),
		.sram(mux_tree_tapbuf_size17_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_1_sram_inv[0:4]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size17 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[44], chanx_left_in[93], chanx_left_in[142], chanx_left_in[191]}),
		.sram(mux_tree_tapbuf_size17_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_2_sram_inv[0:4]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size17 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[43], chanx_left_in[92], chanx_left_in[141], chanx_left_in[190]}),
		.sram(mux_tree_tapbuf_size17_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_3_sram_inv[0:4]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size17 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[42], chanx_left_in[91], chanx_left_in[140], chanx_left_in[189]}),
		.sram(mux_tree_tapbuf_size17_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_4_sram_inv[0:4]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size17 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[41], chanx_left_in[90], chanx_left_in[139], chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size17_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_5_sram_inv[0:4]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size17 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[36], chanx_left_in[85], chanx_left_in[134], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size17_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_6_sram_inv[0:4]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size17 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[35], chanx_left_in[84], chanx_left_in[133], chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size17_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_7_sram_inv[0:4]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size17 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[34], chanx_left_in[83], chanx_left_in[132], chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size17_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_8_sram_inv[0:4]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size17 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[27], chanx_left_in[76], chanx_left_in[125], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size17_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_9_sram_inv[0:4]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size17 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[26], chanx_left_in[75], chanx_left_in[124], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size17_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_10_sram_inv[0:4]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size17 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[24], chanx_left_in[73], chanx_left_in[122], chanx_left_in[171]}),
		.sram(mux_tree_tapbuf_size17_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_11_sram_inv[0:4]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size17 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[17], chanx_left_in[66], chanx_left_in[115], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size17_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_12_sram_inv[0:4]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size17 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[16], chanx_left_in[65], chanx_left_in[114], chanx_left_in[163]}),
		.sram(mux_tree_tapbuf_size17_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_13_sram_inv[0:4]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size17 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[9], chanx_left_in[58], chanx_left_in[107], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size17_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_14_sram_inv[0:4]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size17 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[8], chanx_left_in[57], chanx_left_in[106], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size17_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_15_sram_inv[0:4]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size17 mux_top_track_352 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[5], chanx_left_in[54], chanx_left_in[103], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size17_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_16_sram_inv[0:4]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size17 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[4], chanx_left_in[53], chanx_left_in[102], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size17_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_17_sram_inv[0:4]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size17_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_0_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_1_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_2_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_3_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_4_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_5_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_6_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_7_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_8_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_9_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_10_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_11_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_12_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_13_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_14_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_15_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_16_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_17_sram_inv[0:4]));

	mux_tree_tapbuf_size15 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[48], chanx_left_in[97], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size15_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_0_sram_inv[0:3]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size15 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[47], chanx_left_in[96], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size15_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_1_sram_inv[0:3]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size15 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[46], chanx_left_in[95], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size15_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_2_sram_inv[0:3]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size15_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_0_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_1_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_2_sram_inv[0:3]));

	mux_tree_tapbuf_size16 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[40], chanx_left_in[89], chanx_left_in[138], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size16_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_0_sram_inv[0:4]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size16 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[39], chanx_left_in[88], chanx_left_in[137], chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size16_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_1_sram_inv[0:4]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size16 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[38], chanx_left_in[87], chanx_left_in[136], chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size16_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_2_sram_inv[0:4]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size16 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[37], chanx_left_in[86], chanx_left_in[135], chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size16_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_3_sram_inv[0:4]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size16 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[32], chanx_left_in[81], chanx_left_in[130], chanx_left_in[179]}),
		.sram(mux_tree_tapbuf_size16_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_4_sram_inv[0:4]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size16 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[31], chanx_left_in[80], chanx_left_in[129], chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size16_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_5_sram_inv[0:4]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size16 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[30], chanx_left_in[79], chanx_left_in[128], chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size16_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_6_sram_inv[0:4]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size16 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[29], chanx_left_in[78], chanx_left_in[127], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size16_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_7_sram_inv[0:4]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size16 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[28], chanx_left_in[77], chanx_left_in[126], chanx_left_in[175]}),
		.sram(mux_tree_tapbuf_size16_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_8_sram_inv[0:4]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size16 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[23], chanx_left_in[72], chanx_left_in[121], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size16_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_9_sram_inv[0:4]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size16 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[22], chanx_left_in[71], chanx_left_in[120], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size16_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_10_sram_inv[0:4]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size16 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[21], chanx_left_in[70], chanx_left_in[119], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size16_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_11_sram_inv[0:4]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size16 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[20], chanx_left_in[69], chanx_left_in[118], chanx_left_in[167]}),
		.sram(mux_tree_tapbuf_size16_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_12_sram_inv[0:4]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size16 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[19], chanx_left_in[68], chanx_left_in[117], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size16_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_13_sram_inv[0:4]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size16 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[18], chanx_left_in[67], chanx_left_in[116], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size16_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_14_sram_inv[0:4]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size16 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[15], chanx_left_in[64], chanx_left_in[113], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size16_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_15_sram_inv[0:4]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size16 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[14], chanx_left_in[63], chanx_left_in[112], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size16_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_16_sram_inv[0:4]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size16 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[13], chanx_left_in[62], chanx_left_in[111], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size16_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_17_sram_inv[0:4]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size16 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[12], chanx_left_in[61], chanx_left_in[110], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size16_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_18_sram_inv[0:4]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size16 mux_top_track_304 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[11], chanx_left_in[60], chanx_left_in[109], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size16_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_19_sram_inv[0:4]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size16 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[10], chanx_left_in[59], chanx_left_in[108], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size16_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_20_sram_inv[0:4]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size16 mux_top_track_336 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[7], chanx_left_in[56], chanx_left_in[105], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size16_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_21_sram_inv[0:4]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size16 mux_top_track_344 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[6], chanx_left_in[55], chanx_left_in[104], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size16_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_22_sram_inv[0:4]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size16 mux_top_track_368 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[3], chanx_left_in[52], chanx_left_in[101], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size16_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_23_sram_inv[0:4]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size16 mux_top_track_376 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[2], chanx_left_in[51], chanx_left_in[100], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size16_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_24_sram_inv[0:4]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size16 mux_top_track_384 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[1], chanx_left_in[50], chanx_left_in[99], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size16_25_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_25_sram_inv[0:4]),
		.out(chany_top_out[192]));

	mux_tree_tapbuf_size16_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_0_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_1_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_2_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_3_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_4_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_5_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_6_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_7_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_8_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_9_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_10_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_11_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_12_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_13_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_14_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_15_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_16_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_17_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_18_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_19_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_20_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_21_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_22_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_23_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_24_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_25_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_25_sram_inv[0:4]));

	mux_tree_tapbuf_size18 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[33], chanx_left_in[82], chanx_left_in[131], chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size18_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_0_sram_inv[0:4]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size18 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[25], chanx_left_in[74], chanx_left_in[123], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size18_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_1_sram_inv[0:4]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size18_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_0_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_1_sram_inv[0:4]));

	mux_tree_tapbuf_size6 mux_bottom_track_1 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[1], chanx_left_in[50], chanx_left_in[99], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size6 mux_bottom_track_9 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[2], chanx_left_in[51], chanx_left_in[100], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size6 mux_bottom_track_17 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[3], chanx_left_in[52], chanx_left_in[101], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size6 mux_bottom_track_25 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[4], chanx_left_in[53], chanx_left_in[102], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size6 mux_bottom_track_41 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[6], chanx_left_in[55], chanx_left_in[104], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size6 mux_bottom_track_49 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[7], chanx_left_in[56], chanx_left_in[105], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size6 mux_bottom_track_65 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[9], chanx_left_in[58], chanx_left_in[107], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size6 mux_bottom_track_137 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[18], chanx_left_in[67], chanx_left_in[116], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size6 mux_bottom_track_209 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[27], chanx_left_in[76], chanx_left_in[125], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size6 mux_bottom_track_281 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[36], chanx_left_in[85], chanx_left_in[134], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_9_sram_inv[0:2]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size6 mux_bottom_track_353 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[45], chanx_left_in[94], chanx_left_in[143], chanx_left_in[192]}),
		.sram(mux_tree_tapbuf_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_10_sram_inv[0:2]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_size7 mux_bottom_track_33 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[5], chanx_left_in[54], chanx_left_in[103], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_bottom_track_57 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[8], chanx_left_in[57], chanx_left_in[106], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size5 mux_bottom_track_73 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[10], chanx_left_in[59], chanx_left_in[108], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size5 mux_bottom_track_81 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[11], chanx_left_in[60], chanx_left_in[109], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size5 mux_bottom_track_89 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[12], chanx_left_in[61], chanx_left_in[110], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size5 mux_bottom_track_97 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[13], chanx_left_in[62], chanx_left_in[111], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size5 mux_bottom_track_105 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[14], chanx_left_in[63], chanx_left_in[112], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size5 mux_bottom_track_113 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[15], chanx_left_in[64], chanx_left_in[113], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size5 mux_bottom_track_121 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[16], chanx_left_in[65], chanx_left_in[114], chanx_left_in[163]}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size5 mux_bottom_track_129 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[17], chanx_left_in[66], chanx_left_in[115], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size5 mux_bottom_track_145 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[19], chanx_left_in[68], chanx_left_in[117], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size5 mux_bottom_track_153 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[20], chanx_left_in[69], chanx_left_in[118], chanx_left_in[167]}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size5 mux_bottom_track_161 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[21], chanx_left_in[70], chanx_left_in[119], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size5 mux_bottom_track_169 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[22], chanx_left_in[71], chanx_left_in[120], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size5 mux_bottom_track_177 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[23], chanx_left_in[72], chanx_left_in[121], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size5 mux_bottom_track_185 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[24], chanx_left_in[73], chanx_left_in[122], chanx_left_in[171]}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size5 mux_bottom_track_193 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[25], chanx_left_in[74], chanx_left_in[123], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size5 mux_bottom_track_201 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[26], chanx_left_in[75], chanx_left_in[124], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size5 mux_bottom_track_217 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[28], chanx_left_in[77], chanx_left_in[126], chanx_left_in[175]}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size5 mux_bottom_track_225 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[29], chanx_left_in[78], chanx_left_in[127], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size5 mux_bottom_track_233 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[30], chanx_left_in[79], chanx_left_in[128], chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size5 mux_bottom_track_241 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[31], chanx_left_in[80], chanx_left_in[129], chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size5 mux_bottom_track_249 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[32], chanx_left_in[81], chanx_left_in[130], chanx_left_in[179]}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size5 mux_bottom_track_257 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[33], chanx_left_in[82], chanx_left_in[131], chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size5 mux_bottom_track_265 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[34], chanx_left_in[83], chanx_left_in[132], chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size5 mux_bottom_track_273 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[35], chanx_left_in[84], chanx_left_in[133], chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size5 mux_bottom_track_289 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[37], chanx_left_in[86], chanx_left_in[135], chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size5 mux_bottom_track_297 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[38], chanx_left_in[87], chanx_left_in[136], chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size5 mux_bottom_track_305 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[39], chanx_left_in[88], chanx_left_in[137], chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size5 mux_bottom_track_313 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[40], chanx_left_in[89], chanx_left_in[138], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size5 mux_bottom_track_321 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[41], chanx_left_in[90], chanx_left_in[139], chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size5_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_29_sram_inv[0:2]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size5 mux_bottom_track_329 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[42], chanx_left_in[91], chanx_left_in[140], chanx_left_in[189]}),
		.sram(mux_tree_tapbuf_size5_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_30_sram_inv[0:2]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size5 mux_bottom_track_337 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[43], chanx_left_in[92], chanx_left_in[141], chanx_left_in[190]}),
		.sram(mux_tree_tapbuf_size5_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_31_sram_inv[0:2]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size5 mux_bottom_track_345 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[44], chanx_left_in[93], chanx_left_in[142], chanx_left_in[191]}),
		.sram(mux_tree_tapbuf_size5_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_32_sram_inv[0:2]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size5 mux_bottom_track_385 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[0], chanx_left_in[49], chanx_left_in[98], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size5_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_33_sram_inv[0:2]),
		.out(chany_bottom_out[192]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_29_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_30_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_31_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_32_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_33_sram_inv[0:2]));

	mux_tree_tapbuf_size4 mux_bottom_track_361 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[46], chanx_left_in[95], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size4 mux_bottom_track_369 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[47], chanx_left_in[96], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size4 mux_bottom_track_377 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[48], chanx_left_in[97], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size13 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_0_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size13 mux_left_track_7 (
		.in({chany_bottom_in[2], chany_bottom_in[11], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_1_sram_inv[0:3]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_size13 mux_left_track_19 (
		.in({chany_bottom_in[10], chany_bottom_in[35], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_2_sram_inv[0:3]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_size13 mux_left_track_37 (
		.in({chany_bottom_in[22], chany_bottom_in[71], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_3_sram_inv[0:3]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_size13 mux_left_track_55 (
		.in({chany_bottom_in[34], chany_bottom_in[107], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_4_sram_inv[0:3]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_size13 mux_left_track_73 (
		.in({chany_bottom_in[46], chany_bottom_in[143], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_5_sram_inv[0:3]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size13 mux_left_track_91 (
		.in({chany_bottom_in[58], chany_bottom_in[179], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_6_sram_inv[0:3]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_size13 mux_left_track_109 (
		.in({chany_top_in[185], chany_bottom_in[70], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_7_sram_inv[0:3]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_size13 mux_left_track_127 (
		.in({chany_top_in[173], chany_bottom_in[82], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_8_sram_inv[0:3]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_size13 mux_left_track_163 (
		.in({chany_top_in[149], chany_bottom_in[106], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_9_sram_inv[0:3]),
		.out(chanx_left_out[81]));

	mux_tree_tapbuf_size13 mux_left_track_297 (
		.in({chany_top_in[60], chany_top_in[183], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size13_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_10_sram_inv[0:3]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size13 mux_left_track_315 (
		.in({chany_top_in[48], chany_top_in[147], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size13_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_11_sram_inv[0:3]),
		.out(chanx_left_out[157]));

	mux_tree_tapbuf_size13 mux_left_track_333 (
		.in({chany_top_in[36], chany_top_in[111], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size13_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_12_sram_inv[0:3]),
		.out(chanx_left_out[166]));

	mux_tree_tapbuf_size13_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_163 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_9_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_10_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_315 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_11_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_left_track_333 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_12_sram_inv[0:3]));

	mux_tree_tapbuf_size12 mux_left_track_3 (
		.in({chany_bottom_in[0], chany_bottom_in[3], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_0_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_size12 mux_left_track_9 (
		.in({chany_bottom_in[4], chany_bottom_in[15], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_1_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size12 mux_left_track_11 (
		.in({chany_bottom_in[5], chany_bottom_in[19], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_2_sram_inv[0:3]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_size12 mux_left_track_21 (
		.in({chany_bottom_in[12], chany_bottom_in[39], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_3_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_size12 mux_left_track_23 (
		.in({chany_bottom_in[13], chany_bottom_in[43], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_4_sram_inv[0:3]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_size12 mux_left_track_27 (
		.in({chany_bottom_in[16], chany_bottom_in[51], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_5_sram_inv[0:3]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_size12 mux_left_track_29 (
		.in({chany_bottom_in[17], chany_bottom_in[55], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_6_sram_inv[0:3]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_size12 mux_left_track_31 (
		.in({chany_bottom_in[18], chany_bottom_in[59], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_7_sram_inv[0:3]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_size12 mux_left_track_39 (
		.in({chany_bottom_in[24], chany_bottom_in[75], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_8_sram_inv[0:3]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_size12 mux_left_track_41 (
		.in({chany_bottom_in[25], chany_bottom_in[79], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_9_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size12 mux_left_track_43 (
		.in({chany_bottom_in[26], chany_bottom_in[83], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_10_sram_inv[0:3]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_size12 mux_left_track_47 (
		.in({chany_bottom_in[29], chany_bottom_in[91], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_11_sram_inv[0:3]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_size12 mux_left_track_49 (
		.in({chany_bottom_in[30], chany_bottom_in[95], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_12_sram_inv[0:3]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size12 mux_left_track_51 (
		.in({chany_bottom_in[32], chany_bottom_in[99], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_13_sram_inv[0:3]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_size12 mux_left_track_57 (
		.in({chany_bottom_in[36], chany_bottom_in[111], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_14_sram_inv[0:3]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size12 mux_left_track_59 (
		.in({chany_bottom_in[37], chany_bottom_in[115], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_15_sram_inv[0:3]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_size12 mux_left_track_61 (
		.in({chany_bottom_in[38], chany_bottom_in[119], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_16_sram_inv[0:3]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_size12 mux_left_track_63 (
		.in({chany_bottom_in[40], chany_bottom_in[123], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_17_sram_inv[0:3]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_size12 mux_left_track_67 (
		.in({chany_bottom_in[42], chany_bottom_in[131], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_18_sram_inv[0:3]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_size12 mux_left_track_69 (
		.in({chany_bottom_in[44], chany_bottom_in[135], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_19_sram_inv[0:3]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_size12 mux_left_track_75 (
		.in({chany_bottom_in[48], chany_bottom_in[147], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size12_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_20_sram_inv[0:3]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_size12 mux_left_track_77 (
		.in({chany_bottom_in[49], chany_bottom_in[151], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_21_sram_inv[0:3]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_size12 mux_left_track_79 (
		.in({chany_bottom_in[50], chany_bottom_in[155], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_22_sram_inv[0:3]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_size12 mux_left_track_81 (
		.in({chany_bottom_in[52], chany_bottom_in[159], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_23_sram_inv[0:3]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size12 mux_left_track_83 (
		.in({chany_bottom_in[53], chany_bottom_in[163], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_24_sram_inv[0:3]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_size12 mux_left_track_87 (
		.in({chany_bottom_in[56], chany_bottom_in[171], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_25_sram_inv[0:3]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_size12 mux_left_track_93 (
		.in({chany_bottom_in[60], chany_bottom_in[183], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size12_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_26_sram_inv[0:3]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_size12 mux_left_track_95 (
		.in({chany_bottom_in[61], chany_bottom_in[187], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size12_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_27_sram_inv[0:3]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_size12 mux_left_track_97 (
		.in({chany_bottom_in[62], chany_bottom_in[191], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_28_sram_inv[0:3]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size12 mux_left_track_99 (
		.in({chany_bottom_in[64], chany_bottom_in[192], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_29_sram_inv[0:3]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_size12 mux_left_track_101 (
		.in({chany_top_in[190], chany_bottom_in[65], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_30_sram_inv[0:3]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_size12 mux_left_track_103 (
		.in({chany_top_in[189], chany_bottom_in[66], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_31_sram_inv[0:3]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_size12 mux_left_track_111 (
		.in({chany_top_in[184], chany_bottom_in[72], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_32_sram_inv[0:3]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_size12 mux_left_track_113 (
		.in({chany_top_in[182], chany_bottom_in[73], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size12_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_33_sram_inv[0:3]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size12 mux_left_track_115 (
		.in({chany_top_in[181], chany_bottom_in[74], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size12_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_34_sram_inv[0:3]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_size12 mux_left_track_117 (
		.in({chany_top_in[180], chany_bottom_in[76], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_35_sram_inv[0:3]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_size12 mux_left_track_119 (
		.in({chany_top_in[178], chany_bottom_in[77], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_36_sram_inv[0:3]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_size12 mux_left_track_121 (
		.in({chany_top_in[177], chany_bottom_in[78], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_37_sram_inv[0:3]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size12 mux_left_track_123 (
		.in({chany_top_in[176], chany_bottom_in[80], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_38_sram_inv[0:3]),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_size12 mux_left_track_129 (
		.in({chany_top_in[172], chany_bottom_in[84], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_39_sram_inv[0:3]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size12 mux_left_track_131 (
		.in({chany_top_in[170], chany_bottom_in[85], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_40_sram_inv[0:3]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_size12 mux_left_track_133 (
		.in({chany_top_in[169], chany_bottom_in[86], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size12_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_41_sram_inv[0:3]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_size12 mux_left_track_135 (
		.in({chany_top_in[168], chany_bottom_in[88], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size12_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_42_sram_inv[0:3]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_size12 mux_left_track_137 (
		.in({chany_top_in[166], chany_bottom_in[89], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_43_sram_inv[0:3]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size12 mux_left_track_139 (
		.in({chany_top_in[165], chany_bottom_in[90], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_44_sram_inv[0:3]),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_size12 mux_left_track_141 (
		.in({chany_top_in[164], chany_bottom_in[92], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_45_sram_inv[0:3]),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_size12 mux_left_track_145 (
		.in({chany_top_in[161], chany_bottom_in[94], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_46_sram_inv[0:3]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size12 mux_left_track_147 (
		.in({chany_top_in[160], chany_bottom_in[96], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_47_sram_inv[0:3]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_size12 mux_left_track_149 (
		.in({chany_top_in[158], chany_bottom_in[97], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_48_sram_inv[0:3]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_size12 mux_left_track_151 (
		.in({chany_top_in[157], chany_bottom_in[98], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_49_sram_inv[0:3]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_size12 mux_left_track_153 (
		.in({chany_top_in[156], chany_bottom_in[100], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size12_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_50_sram_inv[0:3]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size12 mux_left_track_155 (
		.in({chany_top_in[154], chany_bottom_in[101], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size12_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_51_sram_inv[0:3]),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_size12 mux_left_track_157 (
		.in({chany_top_in[153], chany_bottom_in[102], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_52_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_52_sram_inv[0:3]),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_size12 mux_left_track_159 (
		.in({chany_top_in[152], chany_bottom_in[104], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_53_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_53_sram_inv[0:3]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_size12 mux_left_track_167 (
		.in({chany_top_in[146], chany_bottom_in[109], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_54_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_54_sram_inv[0:3]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_size12 mux_left_track_169 (
		.in({chany_top_in[145], chany_bottom_in[110], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_55_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_55_sram_inv[0:3]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size12 mux_left_track_171 (
		.in({chany_top_in[144], chany_bottom_in[112], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_56_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_56_sram_inv[0:3]),
		.out(chanx_left_out[85]));

	mux_tree_tapbuf_size12 mux_left_track_173 (
		.in({chany_top_in[142], chany_bottom_in[113], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_57_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_57_sram_inv[0:3]),
		.out(chanx_left_out[86]));

	mux_tree_tapbuf_size12 mux_left_track_175 (
		.in({chany_top_in[141], chany_bottom_in[114], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_58_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_58_sram_inv[0:3]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_size12 mux_left_track_177 (
		.in({chany_top_in[140], chany_bottom_in[116], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_59_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_59_sram_inv[0:3]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size12 mux_left_track_189 (
		.in({chany_top_in[132], chany_bottom_in[124], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_60_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_60_sram_inv[0:3]),
		.out(chanx_left_out[94]));

	mux_tree_tapbuf_size12 mux_left_track_193 (
		.in({chany_top_in[129], chany_bottom_in[126], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_61_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_61_sram_inv[0:3]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size12 mux_left_track_195 (
		.in({chany_top_in[128], chany_bottom_in[128], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_62_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_62_sram_inv[0:3]),
		.out(chanx_left_out[97]));

	mux_tree_tapbuf_size12 mux_left_track_207 (
		.in({chany_top_in[120], chany_bottom_in[136], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_63_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_63_sram_inv[0:3]),
		.out(chanx_left_out[103]));

	mux_tree_tapbuf_size12 mux_left_track_213 (
		.in({chany_top_in[116], chany_bottom_in[140], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_64_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_64_sram_inv[0:3]),
		.out(chanx_left_out[106]));

	mux_tree_tapbuf_size12 mux_left_track_217 (
		.in({chany_top_in[113], chany_bottom_in[142], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_65_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_65_sram_inv[0:3]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size12 mux_left_track_225 (
		.in({chany_top_in[108], chany_bottom_in[148], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_66_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_66_sram_inv[0:3]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size12 mux_left_track_235 (
		.in({chany_top_in[101], chany_bottom_in[154], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_67_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_67_sram_inv[0:3]),
		.out(chanx_left_out[117]));

	mux_tree_tapbuf_size12 mux_left_track_237 (
		.in({chany_top_in[100], chany_bottom_in[156], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_68_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_68_sram_inv[0:3]),
		.out(chanx_left_out[118]));

	mux_tree_tapbuf_size12 mux_left_track_243 (
		.in({chany_top_in[96], chany_bottom_in[160], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_69_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_69_sram_inv[0:3]),
		.out(chanx_left_out[121]));

	mux_tree_tapbuf_size12 mux_left_track_253 (
		.in({chany_top_in[89], chany_bottom_in[166], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_70_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_70_sram_inv[0:3]),
		.out(chanx_left_out[126]));

	mux_tree_tapbuf_size12 mux_left_track_255 (
		.in({chany_top_in[88], chany_bottom_in[168], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_71_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_71_sram_inv[0:3]),
		.out(chanx_left_out[127]));

	mux_tree_tapbuf_size12 mux_left_track_257 (
		.in({chany_top_in[86], chany_bottom_in[169], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_72_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_72_sram_inv[0:3]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size12 mux_left_track_261 (
		.in({chany_top_in[84], chany_bottom_in[172], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_73_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_73_sram_inv[0:3]),
		.out(chanx_left_out[130]));

	mux_tree_tapbuf_size12 mux_left_track_273 (
		.in({chany_top_in[76], chany_bottom_in[180], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_74_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_74_sram_inv[0:3]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size12 mux_left_track_275 (
		.in({chany_top_in[74], chany_bottom_in[181], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_75_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_75_sram_inv[0:3]),
		.out(chanx_left_out[137]));

	mux_tree_tapbuf_size12 mux_left_track_277 (
		.in({chany_top_in[73], chany_bottom_in[182], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_76_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_76_sram_inv[0:3]),
		.out(chanx_left_out[138]));

	mux_tree_tapbuf_size12 mux_left_track_279 (
		.in({chany_top_in[72], chany_bottom_in[184], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_77_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_77_sram_inv[0:3]),
		.out(chanx_left_out[139]));

	mux_tree_tapbuf_size12 mux_left_track_293 (
		.in({chany_top_in[62], chany_top_in[191], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_78_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_78_sram_inv[0:3]),
		.out(chanx_left_out[146]));

	mux_tree_tapbuf_size12 mux_left_track_295 (
		.in({chany_top_in[61], chany_top_in[187], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_79_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_79_sram_inv[0:3]),
		.out(chanx_left_out[147]));

	mux_tree_tapbuf_size12 mux_left_track_313 (
		.in({chany_top_in[49], chany_top_in[151], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_80_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_80_sram_inv[0:3]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size12 mux_left_track_317 (
		.in({chany_top_in[46], chany_top_in[143], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_81_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_81_sram_inv[0:3]),
		.out(chanx_left_out[158]));

	mux_tree_tapbuf_size12 mux_left_track_335 (
		.in({chany_top_in[34], chany_top_in[107], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_82_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_82_sram_inv[0:3]),
		.out(chanx_left_out[167]));

	mux_tree_tapbuf_size12 mux_left_track_337 (
		.in({chany_top_in[33], chany_top_in[103], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_83_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_83_sram_inv[0:3]),
		.out(chanx_left_out[168]));

	mux_tree_tapbuf_size12 mux_left_track_353 (
		.in({chany_top_in[22], chany_top_in[71], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_84_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_84_sram_inv[0:3]),
		.out(chanx_left_out[176]));

	mux_tree_tapbuf_size12 mux_left_track_355 (
		.in({chany_top_in[21], chany_top_in[67], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_85_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_85_sram_inv[0:3]),
		.out(chanx_left_out[177]));

	mux_tree_tapbuf_size12 mux_left_track_357 (
		.in({chany_top_in[20], chany_top_in[63], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_86_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_86_sram_inv[0:3]),
		.out(chanx_left_out[178]));

	mux_tree_tapbuf_size12 mux_left_track_369 (
		.in({chany_top_in[12], chany_top_in[39], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size12_87_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_87_sram_inv[0:3]),
		.out(chanx_left_out[184]));

	mux_tree_tapbuf_size12 mux_left_track_373 (
		.in({chany_top_in[9], chany_top_in[31], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_88_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_88_sram_inv[0:3]),
		.out(chanx_left_out[186]));

	mux_tree_tapbuf_size12 mux_left_track_375 (
		.in({chany_top_in[8], chany_top_in[27], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_89_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_89_sram_inv[0:3]),
		.out(chanx_left_out[187]));

	mux_tree_tapbuf_size12_mem mem_left_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_16_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_17_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_18_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_19_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_20_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_21_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_22_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_23_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_24_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_25_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_26_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_27_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_28_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_29_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_30_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_31_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_32_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_33_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_34_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_35_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_36_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_37_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_38_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_39_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_40_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_41_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_42_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_43_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_44_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_45_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_46_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_147 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_47_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_149 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_48_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_151 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_49_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_50_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_155 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_51_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_157 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_52_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_52_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_159 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_53_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_53_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_167 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_54_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_54_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_55_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_55_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_171 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_56_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_56_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_173 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_57_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_57_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_175 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_58_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_58_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_59_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_59_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_189 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_60_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_60_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_61_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_61_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_195 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_62_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_62_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_207 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_63_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_63_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_213 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_64_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_64_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_65_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_65_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_66_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_66_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_235 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_67_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_67_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_237 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_68_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_68_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_243 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_69_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_69_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_253 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_70_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_70_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_255 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_71_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_71_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_72_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_72_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_261 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_73_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_73_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_74_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_74_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_275 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_75_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_75_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_277 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_76_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_76_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_279 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_77_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_77_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_293 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_78_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_78_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_295 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_79_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_79_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_80_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_80_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_317 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_81_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_81_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_335 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_82_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_82_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_83_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_83_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_84_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_84_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_355 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_85_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_85_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_357 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_86_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_86_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_87_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_87_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_373 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_88_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_88_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_375 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_89_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_89_sram_inv[0:3]));

	mux_tree_tapbuf_size11 mux_left_track_5 (
		.in({chany_bottom_in[1], chany_bottom_in[7], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_0_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_size11 mux_left_track_13 (
		.in({chany_bottom_in[6], chany_bottom_in[23], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_1_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_size11 mux_left_track_15 (
		.in({chany_bottom_in[8], chany_bottom_in[27], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_2_sram_inv[0:3]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_size11 mux_left_track_17 (
		.in({chany_bottom_in[9], chany_bottom_in[31], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_3_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size11 mux_left_track_25 (
		.in({chany_bottom_in[14], chany_bottom_in[47], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_4_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size11 mux_left_track_33 (
		.in({chany_bottom_in[20], chany_bottom_in[63], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_5_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size11 mux_left_track_35 (
		.in({chany_bottom_in[21], chany_bottom_in[67], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_6_sram_inv[0:3]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_size11 mux_left_track_53 (
		.in({chany_bottom_in[33], chany_bottom_in[103], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_7_sram_inv[0:3]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_size11 mux_left_track_65 (
		.in({chany_bottom_in[41], chany_bottom_in[127], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_8_sram_inv[0:3]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size11 mux_left_track_71 (
		.in({chany_bottom_in[45], chany_bottom_in[139], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_9_sram_inv[0:3]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_size11 mux_left_track_85 (
		.in({chany_bottom_in[54], chany_bottom_in[167], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_10_sram_inv[0:3]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_size11 mux_left_track_89 (
		.in({chany_bottom_in[57], chany_bottom_in[175], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_11_sram_inv[0:3]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size11 mux_left_track_105 (
		.in({chany_top_in[188], chany_bottom_in[68], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_12_sram_inv[0:3]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size11 mux_left_track_107 (
		.in({chany_top_in[186], chany_bottom_in[69], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size11_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_13_sram_inv[0:3]),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_size11 mux_left_track_143 (
		.in({chany_top_in[162], chany_bottom_in[93], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_14_sram_inv[0:3]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_size11 mux_left_track_161 (
		.in({chany_top_in[150], chany_bottom_in[105], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_15_sram_inv[0:3]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size11 mux_left_track_165 (
		.in({chany_top_in[148], chany_bottom_in[108], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_16_sram_inv[0:3]),
		.out(chanx_left_out[82]));

	mux_tree_tapbuf_size11 mux_left_track_181 (
		.in({chany_top_in[137], chany_bottom_in[118], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_17_sram_inv[0:3]),
		.out(chanx_left_out[90]));

	mux_tree_tapbuf_size11 mux_left_track_183 (
		.in({chany_top_in[136], chany_bottom_in[120], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_18_sram_inv[0:3]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_size11 mux_left_track_185 (
		.in({chany_top_in[134], chany_bottom_in[121], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_19_sram_inv[0:3]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size11 mux_left_track_187 (
		.in({chany_top_in[133], chany_bottom_in[122], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_20_sram_inv[0:3]),
		.out(chanx_left_out[93]));

	mux_tree_tapbuf_size11 mux_left_track_197 (
		.in({chany_top_in[126], chany_bottom_in[129], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size11_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_21_sram_inv[0:3]),
		.out(chanx_left_out[98]));

	mux_tree_tapbuf_size11 mux_left_track_199 (
		.in({chany_top_in[125], chany_bottom_in[130], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_22_sram_inv[0:3]),
		.out(chanx_left_out[99]));

	mux_tree_tapbuf_size11 mux_left_track_201 (
		.in({chany_top_in[124], chany_bottom_in[132], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_23_sram_inv[0:3]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size11 mux_left_track_203 (
		.in({chany_top_in[122], chany_bottom_in[133], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_24_sram_inv[0:3]),
		.out(chanx_left_out[101]));

	mux_tree_tapbuf_size11 mux_left_track_205 (
		.in({chany_top_in[121], chany_bottom_in[134], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_25_sram_inv[0:3]),
		.out(chanx_left_out[102]));

	mux_tree_tapbuf_size11 mux_left_track_209 (
		.in({chany_top_in[118], chany_bottom_in[137], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_26_sram_inv[0:3]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size11 mux_left_track_215 (
		.in({chany_top_in[114], chany_bottom_in[141], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size11_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_27_sram_inv[0:3]),
		.out(chanx_left_out[107]));

	mux_tree_tapbuf_size11 mux_left_track_219 (
		.in({chany_top_in[112], chany_bottom_in[144], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_28_sram_inv[0:3]),
		.out(chanx_left_out[109]));

	mux_tree_tapbuf_size11 mux_left_track_221 (
		.in({chany_top_in[110], chany_bottom_in[145], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_29_sram_inv[0:3]),
		.out(chanx_left_out[110]));

	mux_tree_tapbuf_size11 mux_left_track_223 (
		.in({chany_top_in[109], chany_bottom_in[146], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_30_sram_inv[0:3]),
		.out(chanx_left_out[111]));

	mux_tree_tapbuf_size11 mux_left_track_227 (
		.in({chany_top_in[106], chany_bottom_in[149], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_31_sram_inv[0:3]),
		.out(chanx_left_out[113]));

	mux_tree_tapbuf_size11 mux_left_track_229 (
		.in({chany_top_in[105], chany_bottom_in[150], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_32_sram_inv[0:3]),
		.out(chanx_left_out[114]));

	mux_tree_tapbuf_size11 mux_left_track_233 (
		.in({chany_top_in[102], chany_bottom_in[153], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size11_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_33_sram_inv[0:3]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size11 mux_left_track_239 (
		.in({chany_top_in[98], chany_bottom_in[157], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_34_sram_inv[0:3]),
		.out(chanx_left_out[119]));

	mux_tree_tapbuf_size11 mux_left_track_241 (
		.in({chany_top_in[97], chany_bottom_in[158], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_35_sram_inv[0:3]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size11 mux_left_track_245 (
		.in({chany_top_in[94], chany_bottom_in[161], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_36_sram_inv[0:3]),
		.out(chanx_left_out[122]));

	mux_tree_tapbuf_size11 mux_left_track_247 (
		.in({chany_top_in[93], chany_bottom_in[162], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_37_sram_inv[0:3]),
		.out(chanx_left_out[123]));

	mux_tree_tapbuf_size11 mux_left_track_249 (
		.in({chany_top_in[92], chany_bottom_in[164], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_38_sram_inv[0:3]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size11 mux_left_track_259 (
		.in({chany_top_in[85], chany_bottom_in[170], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_39_sram_inv[0:3]),
		.out(chanx_left_out[129]));

	mux_tree_tapbuf_size11 mux_left_track_263 (
		.in({chany_top_in[82], chany_bottom_in[173], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_40_sram_inv[0:3]),
		.out(chanx_left_out[131]));

	mux_tree_tapbuf_size11 mux_left_track_265 (
		.in({chany_top_in[81], chany_bottom_in[174], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_41_sram_inv[0:3]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size11 mux_left_track_267 (
		.in({chany_top_in[80], chany_bottom_in[176], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_42_sram_inv[0:3]),
		.out(chanx_left_out[133]));

	mux_tree_tapbuf_size11 mux_left_track_281 (
		.in({chany_top_in[70], chany_bottom_in[185], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_43_sram_inv[0:3]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size11 mux_left_track_283 (
		.in({chany_top_in[69], chany_bottom_in[186], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_44_sram_inv[0:3]),
		.out(chanx_left_out[141]));

	mux_tree_tapbuf_size11 mux_left_track_285 (
		.in({chany_top_in[68], chany_bottom_in[188], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_45_sram_inv[0:3]),
		.out(chanx_left_out[142]));

	mux_tree_tapbuf_size11 mux_left_track_289 (
		.in({chany_top_in[65], chany_bottom_in[190], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_46_sram_inv[0:3]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size11 mux_left_track_299 (
		.in({chany_top_in[58], chany_top_in[179], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_47_sram_inv[0:3]),
		.out(chanx_left_out[149]));

	mux_tree_tapbuf_size11 mux_left_track_301 (
		.in({chany_top_in[57], chany_top_in[175], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_48_sram_inv[0:3]),
		.out(chanx_left_out[150]));

	mux_tree_tapbuf_size11 mux_left_track_303 (
		.in({chany_top_in[56], chany_top_in[171], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_49_sram_inv[0:3]),
		.out(chanx_left_out[151]));

	mux_tree_tapbuf_size11 mux_left_track_307 (
		.in({chany_top_in[53], chany_top_in[163], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_50_sram_inv[0:3]),
		.out(chanx_left_out[153]));

	mux_tree_tapbuf_size11 mux_left_track_309 (
		.in({chany_top_in[52], chany_top_in[159], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_51_sram_inv[0:3]),
		.out(chanx_left_out[154]));

	mux_tree_tapbuf_size11 mux_left_track_319 (
		.in({chany_top_in[45], chany_top_in[139], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_52_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_52_sram_inv[0:3]),
		.out(chanx_left_out[159]));

	mux_tree_tapbuf_size11 mux_left_track_321 (
		.in({chany_top_in[44], chany_top_in[135], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_53_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_53_sram_inv[0:3]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size11 mux_left_track_325 (
		.in({chany_top_in[41], chany_top_in[127], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_54_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_54_sram_inv[0:3]),
		.out(chanx_left_out[162]));

	mux_tree_tapbuf_size11 mux_left_track_327 (
		.in({chany_top_in[40], chany_top_in[123], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_55_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_55_sram_inv[0:3]),
		.out(chanx_left_out[163]));

	mux_tree_tapbuf_size11 mux_left_track_329 (
		.in({chany_top_in[38], chany_top_in[119], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_56_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_56_sram_inv[0:3]),
		.out(chanx_left_out[164]));

	mux_tree_tapbuf_size11 mux_left_track_339 (
		.in({chany_top_in[32], chany_top_in[99], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_57_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_57_sram_inv[0:3]),
		.out(chanx_left_out[169]));

	mux_tree_tapbuf_size11 mux_left_track_343 (
		.in({chany_top_in[29], chany_top_in[91], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_58_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_58_sram_inv[0:3]),
		.out(chanx_left_out[171]));

	mux_tree_tapbuf_size11 mux_left_track_345 (
		.in({chany_top_in[28], chany_top_in[87], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_59_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_59_sram_inv[0:3]),
		.out(chanx_left_out[172]));

	mux_tree_tapbuf_size11 mux_left_track_347 (
		.in({chany_top_in[26], chany_top_in[83], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_60_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_60_sram_inv[0:3]),
		.out(chanx_left_out[173]));

	mux_tree_tapbuf_size11 mux_left_track_349 (
		.in({chany_top_in[25], chany_top_in[79], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size11_61_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_61_sram_inv[0:3]),
		.out(chanx_left_out[174]));

	mux_tree_tapbuf_size11 mux_left_track_351 (
		.in({chany_top_in[24], chany_top_in[75], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size11_62_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_62_sram_inv[0:3]),
		.out(chanx_left_out[175]));

	mux_tree_tapbuf_size11 mux_left_track_361 (
		.in({chany_top_in[17], chany_top_in[55], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_63_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_63_sram_inv[0:3]),
		.out(chanx_left_out[180]));

	mux_tree_tapbuf_size11 mux_left_track_363 (
		.in({chany_top_in[16], chany_top_in[51], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_64_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_64_sram_inv[0:3]),
		.out(chanx_left_out[181]));

	mux_tree_tapbuf_size11 mux_left_track_365 (
		.in({chany_top_in[14], chany_top_in[47], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_65_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_65_sram_inv[0:3]),
		.out(chanx_left_out[182]));

	mux_tree_tapbuf_size11 mux_left_track_367 (
		.in({chany_top_in[13], chany_top_in[43], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size11_66_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_66_sram_inv[0:3]),
		.out(chanx_left_out[183]));

	mux_tree_tapbuf_size11 mux_left_track_377 (
		.in({chany_top_in[6], chany_top_in[23], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size11_67_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_67_sram_inv[0:3]),
		.out(chanx_left_out[188]));

	mux_tree_tapbuf_size11 mux_left_track_379 (
		.in({chany_top_in[5], chany_top_in[19], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_68_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_68_sram_inv[0:3]),
		.out(chanx_left_out[189]));

	mux_tree_tapbuf_size11 mux_left_track_381 (
		.in({chany_top_in[4], chany_top_in[15], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_69_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_69_sram_inv[0:3]),
		.out(chanx_left_out[190]));

	mux_tree_tapbuf_size11 mux_left_track_383 (
		.in({chany_top_in[2], chany_top_in[11], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_70_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_70_sram_inv[0:3]),
		.out(chanx_left_out[191]));

	mux_tree_tapbuf_size11 mux_left_track_385 (
		.in({chany_top_in[1], chany_top_in[7], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size11_71_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_71_sram_inv[0:3]),
		.out(chanx_left_out[192]));

	mux_tree_tapbuf_size11_mem mem_left_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_12_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_13_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_14_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_15_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_165 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_16_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_181 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_17_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_183 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_18_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_19_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_187 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_20_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_197 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_21_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_199 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_22_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_23_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_203 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_24_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_205 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_25_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_26_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_215 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_27_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_219 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_28_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_221 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_29_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_223 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_30_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_227 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_31_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_229 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_32_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_33_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_239 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_34_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_35_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_245 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_36_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_247 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_37_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_38_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_259 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_39_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_263 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_40_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_41_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_267 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_42_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_43_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_283 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_44_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_285 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_45_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_46_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_299 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_47_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_301 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_48_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_303 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_49_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_307 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_50_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_309 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_51_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_319 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_52_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_52_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_53_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_53_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_325 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_54_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_54_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_327 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_55_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_55_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_56_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_56_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_339 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_57_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_57_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_343 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_58_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_58_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_59_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_59_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_347 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_60_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_60_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_349 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_61_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_61_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_351 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_62_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_62_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_63_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_63_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_363 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_64_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_64_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_365 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_65_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_65_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_367 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_66_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_66_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_67_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_67_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_379 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_68_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_68_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_381 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_69_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_69_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_383 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_70_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_70_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_70_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_71_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_71_sram_inv[0:3]));

	mux_tree_tapbuf_size10 mux_left_track_45 (
		.in({chany_bottom_in[28], chany_bottom_in[87], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_0_sram_inv[0:3]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_size10 mux_left_track_125 (
		.in({chany_top_in[174], chany_bottom_in[81], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_1_sram_inv[0:3]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_size10 mux_left_track_179 (
		.in({chany_top_in[138], chany_bottom_in[117], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_2_sram_inv[0:3]),
		.out(chanx_left_out[89]));

	mux_tree_tapbuf_size10 mux_left_track_191 (
		.in({chany_top_in[130], chany_bottom_in[125], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_3_sram_inv[0:3]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_size10 mux_left_track_211 (
		.in({chany_top_in[117], chany_bottom_in[138], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_4_sram_inv[0:3]),
		.out(chanx_left_out[105]));

	mux_tree_tapbuf_size10 mux_left_track_231 (
		.in({chany_top_in[104], chany_bottom_in[152], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_5_sram_inv[0:3]),
		.out(chanx_left_out[115]));

	mux_tree_tapbuf_size10 mux_left_track_269 (
		.in({chany_top_in[78], chany_bottom_in[177], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size10_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_6_sram_inv[0:3]),
		.out(chanx_left_out[134]));

	mux_tree_tapbuf_size10 mux_left_track_271 (
		.in({chany_top_in[77], chany_bottom_in[178], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_7_sram_inv[0:3]),
		.out(chanx_left_out[135]));

	mux_tree_tapbuf_size10 mux_left_track_287 (
		.in({chany_top_in[66], chany_bottom_in[189], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size10_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_8_sram_inv[0:3]),
		.out(chanx_left_out[143]));

	mux_tree_tapbuf_size10 mux_left_track_291 (
		.in({chany_top_in[64], chany_top_in[192], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_9_sram_inv[0:3]),
		.out(chanx_left_out[145]));

	mux_tree_tapbuf_size10 mux_left_track_305 (
		.in({chany_top_in[54], chany_top_in[167], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size10_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_10_sram_inv[0:3]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size10 mux_left_track_311 (
		.in({chany_top_in[50], chany_top_in[155], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_11_sram_inv[0:3]),
		.out(chanx_left_out[155]));

	mux_tree_tapbuf_size10 mux_left_track_323 (
		.in({chany_top_in[42], chany_top_in[131], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size10_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_12_sram_inv[0:3]),
		.out(chanx_left_out[161]));

	mux_tree_tapbuf_size10 mux_left_track_331 (
		.in({chany_top_in[37], chany_top_in[115], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_13_sram_inv[0:3]),
		.out(chanx_left_out[165]));

	mux_tree_tapbuf_size10 mux_left_track_341 (
		.in({chany_top_in[30], chany_top_in[95], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size10_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_14_sram_inv[0:3]),
		.out(chanx_left_out[170]));

	mux_tree_tapbuf_size10 mux_left_track_359 (
		.in({chany_top_in[18], chany_top_in[59], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size10_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_15_sram_inv[0:3]),
		.out(chanx_left_out[179]));

	mux_tree_tapbuf_size10 mux_left_track_371 (
		.in({chany_top_in[10], chany_top_in[35], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_16_sram_inv[0:3]),
		.out(chanx_left_out[185]));

	mux_tree_tapbuf_size10_mem mem_left_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_179 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_191 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_3_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_211 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_4_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_231 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_5_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_269 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_6_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_271 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_7_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_287 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_8_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_291 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_9_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_10_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_311 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_11_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_323 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_12_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_331 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_13_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_341 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_14_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_359 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_15_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_371 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_16_sram_inv[0:3]));

	mux_tree_tapbuf_size9 mux_left_track_251 (
		.in({chany_top_in[90], chany_bottom_in[165], left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_0_sram_inv[0:3]),
		.out(chanx_left_out[125]));

	mux_tree_tapbuf_size9_mem mem_left_track_251 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_0_sram_inv[0:3]));

endmodule
// ----- END Verilog module for sb_4__1_ -----

//----- Default net type -----
`default_nettype wire



