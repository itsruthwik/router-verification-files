//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Connection Blocks[5][6]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul  7 20:54:35 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for cby_5__6_ -----
module cby_5__6_(prog_clk,
                 chany_bottom_in,
                 chany_top_in,
                 ccff_head,
                 chany_bottom_out,
                 chany_top_out,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_0_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_1_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_2_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_3_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_4_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_5_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_6_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_7_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_8_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_9_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_10_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_11_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_12_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_13_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_14_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_15_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_16_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_17_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_18_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_19_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_20_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_21_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_22_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_23_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_24_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_25_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_26_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_27_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_28_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_29_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_30_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_31_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_32_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_33_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_34_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_35_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_36_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_37_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_38_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_39_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_40_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_41_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_42_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_43_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_44_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_45_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_46_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_47_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_48_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_49_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_50_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_51_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_52_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_53_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_54_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_55_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_56_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_57_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_58_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_59_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_60_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_61_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_62_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_63_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_64_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_65_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_66_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_67_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_68_,
                 right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_69_,
                 right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_0_,
                 right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_1_,
                 right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_2_,
                 right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_0_,
                 right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_1_,
                 right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_2_,
                 left_grid_right_width_0_height_0_subtile_0__pin_I_1_,
                 left_grid_right_width_0_height_0_subtile_0__pin_I_5_,
                 left_grid_right_width_0_height_0_subtile_0__pin_I_9_,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:295] chany_bottom_in;
//----- INPUT PORTS -----
input [0:295] chany_top_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:295] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:295] chany_top_out;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_0_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_1_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_2_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_3_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_4_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_5_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_6_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_7_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_8_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_9_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_10_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_11_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_12_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_13_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_14_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_15_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_16_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_17_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_18_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_19_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_20_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_21_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_22_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_23_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_24_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_25_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_26_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_27_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_28_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_29_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_30_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_31_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_32_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_33_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_34_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_35_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_36_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_37_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_38_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_39_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_40_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_41_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_42_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_43_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_44_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_45_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_46_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_47_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_48_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_49_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_50_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_51_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_52_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_53_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_54_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_55_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_56_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_57_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_58_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_59_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_60_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_61_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_62_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_63_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_64_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_65_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_66_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_67_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_68_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_69_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_0_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_1_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_2_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_0_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_1_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_2_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:6] mux_tree_tapbuf_size100_0_sram;
wire [0:6] mux_tree_tapbuf_size100_0_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_10_sram;
wire [0:6] mux_tree_tapbuf_size100_10_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_11_sram;
wire [0:6] mux_tree_tapbuf_size100_11_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_12_sram;
wire [0:6] mux_tree_tapbuf_size100_12_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_13_sram;
wire [0:6] mux_tree_tapbuf_size100_13_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_14_sram;
wire [0:6] mux_tree_tapbuf_size100_14_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_15_sram;
wire [0:6] mux_tree_tapbuf_size100_15_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_16_sram;
wire [0:6] mux_tree_tapbuf_size100_16_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_17_sram;
wire [0:6] mux_tree_tapbuf_size100_17_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_18_sram;
wire [0:6] mux_tree_tapbuf_size100_18_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_19_sram;
wire [0:6] mux_tree_tapbuf_size100_19_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_1_sram;
wire [0:6] mux_tree_tapbuf_size100_1_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_20_sram;
wire [0:6] mux_tree_tapbuf_size100_20_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_21_sram;
wire [0:6] mux_tree_tapbuf_size100_21_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_22_sram;
wire [0:6] mux_tree_tapbuf_size100_22_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_23_sram;
wire [0:6] mux_tree_tapbuf_size100_23_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_24_sram;
wire [0:6] mux_tree_tapbuf_size100_24_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_25_sram;
wire [0:6] mux_tree_tapbuf_size100_25_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_26_sram;
wire [0:6] mux_tree_tapbuf_size100_26_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_27_sram;
wire [0:6] mux_tree_tapbuf_size100_27_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_28_sram;
wire [0:6] mux_tree_tapbuf_size100_28_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_29_sram;
wire [0:6] mux_tree_tapbuf_size100_29_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_2_sram;
wire [0:6] mux_tree_tapbuf_size100_2_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_30_sram;
wire [0:6] mux_tree_tapbuf_size100_30_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_31_sram;
wire [0:6] mux_tree_tapbuf_size100_31_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_32_sram;
wire [0:6] mux_tree_tapbuf_size100_32_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_33_sram;
wire [0:6] mux_tree_tapbuf_size100_33_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_34_sram;
wire [0:6] mux_tree_tapbuf_size100_34_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_35_sram;
wire [0:6] mux_tree_tapbuf_size100_35_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_36_sram;
wire [0:6] mux_tree_tapbuf_size100_36_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_37_sram;
wire [0:6] mux_tree_tapbuf_size100_37_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_38_sram;
wire [0:6] mux_tree_tapbuf_size100_38_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_39_sram;
wire [0:6] mux_tree_tapbuf_size100_39_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_3_sram;
wire [0:6] mux_tree_tapbuf_size100_3_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_40_sram;
wire [0:6] mux_tree_tapbuf_size100_40_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_41_sram;
wire [0:6] mux_tree_tapbuf_size100_41_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_42_sram;
wire [0:6] mux_tree_tapbuf_size100_42_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_43_sram;
wire [0:6] mux_tree_tapbuf_size100_43_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_44_sram;
wire [0:6] mux_tree_tapbuf_size100_44_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_45_sram;
wire [0:6] mux_tree_tapbuf_size100_45_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_46_sram;
wire [0:6] mux_tree_tapbuf_size100_46_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_47_sram;
wire [0:6] mux_tree_tapbuf_size100_47_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_48_sram;
wire [0:6] mux_tree_tapbuf_size100_48_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_49_sram;
wire [0:6] mux_tree_tapbuf_size100_49_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_4_sram;
wire [0:6] mux_tree_tapbuf_size100_4_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_50_sram;
wire [0:6] mux_tree_tapbuf_size100_50_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_51_sram;
wire [0:6] mux_tree_tapbuf_size100_51_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_52_sram;
wire [0:6] mux_tree_tapbuf_size100_52_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_53_sram;
wire [0:6] mux_tree_tapbuf_size100_53_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_54_sram;
wire [0:6] mux_tree_tapbuf_size100_54_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_55_sram;
wire [0:6] mux_tree_tapbuf_size100_55_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_56_sram;
wire [0:6] mux_tree_tapbuf_size100_56_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_57_sram;
wire [0:6] mux_tree_tapbuf_size100_57_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_58_sram;
wire [0:6] mux_tree_tapbuf_size100_58_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_59_sram;
wire [0:6] mux_tree_tapbuf_size100_59_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_5_sram;
wire [0:6] mux_tree_tapbuf_size100_5_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_60_sram;
wire [0:6] mux_tree_tapbuf_size100_60_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_61_sram;
wire [0:6] mux_tree_tapbuf_size100_61_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_62_sram;
wire [0:6] mux_tree_tapbuf_size100_62_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_63_sram;
wire [0:6] mux_tree_tapbuf_size100_63_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_64_sram;
wire [0:6] mux_tree_tapbuf_size100_64_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_65_sram;
wire [0:6] mux_tree_tapbuf_size100_65_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_66_sram;
wire [0:6] mux_tree_tapbuf_size100_66_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_67_sram;
wire [0:6] mux_tree_tapbuf_size100_67_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_68_sram;
wire [0:6] mux_tree_tapbuf_size100_68_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_69_sram;
wire [0:6] mux_tree_tapbuf_size100_69_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_6_sram;
wire [0:6] mux_tree_tapbuf_size100_6_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_70_sram;
wire [0:6] mux_tree_tapbuf_size100_70_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_71_sram;
wire [0:6] mux_tree_tapbuf_size100_71_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_72_sram;
wire [0:6] mux_tree_tapbuf_size100_72_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_73_sram;
wire [0:6] mux_tree_tapbuf_size100_73_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_74_sram;
wire [0:6] mux_tree_tapbuf_size100_74_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_75_sram;
wire [0:6] mux_tree_tapbuf_size100_75_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_76_sram;
wire [0:6] mux_tree_tapbuf_size100_76_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_77_sram;
wire [0:6] mux_tree_tapbuf_size100_77_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_78_sram;
wire [0:6] mux_tree_tapbuf_size100_78_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_7_sram;
wire [0:6] mux_tree_tapbuf_size100_7_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_8_sram;
wire [0:6] mux_tree_tapbuf_size100_8_sram_inv;
wire [0:6] mux_tree_tapbuf_size100_9_sram;
wire [0:6] mux_tree_tapbuf_size100_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size100_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size100_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[0] = chany_bottom_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[4] = chany_bottom_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chany_bottom_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[12] = chany_bottom_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[16] = chany_bottom_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[20] = chany_bottom_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[24] = chany_bottom_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[28] = chany_bottom_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[32] = chany_bottom_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[36] = chany_bottom_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[40] = chany_bottom_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chany_bottom_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[48] = chany_bottom_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[52] = chany_bottom_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[56] = chany_bottom_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chany_bottom_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[64] = chany_bottom_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[66];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[68] = chany_bottom_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[70];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[72] = chany_bottom_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[74];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[76] = chany_bottom_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[78];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chany_bottom_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[82];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[84] = chany_bottom_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[86];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[88] = chany_bottom_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[90];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[92] = chany_bottom_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[94];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[95];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[96] = chany_bottom_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[98];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[100] = chany_bottom_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[102];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[103];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[104] = chany_bottom_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[106];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[107];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[108] = chany_bottom_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[110];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[111];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[112] = chany_bottom_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[114];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[115];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[116] = chany_bottom_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[118];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[119];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[120] = chany_bottom_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[122];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[123];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[124] = chany_bottom_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[126];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[127];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[128] = chany_bottom_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[130];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[131];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[132] = chany_bottom_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[134];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[135];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[136] = chany_bottom_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[138];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[139];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[140] = chany_bottom_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[142];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[143];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[144] = chany_bottom_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[146];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[147];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[148] = chany_bottom_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[150];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[151];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[152] = chany_bottom_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[154];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[155];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[156] = chany_bottom_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[158];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[159];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[160] = chany_bottom_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[162];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[163];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[164] = chany_bottom_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[166];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[167];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[168] = chany_bottom_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[170];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[171];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[172] = chany_bottom_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[174];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[175];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[176] = chany_bottom_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[178];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[179];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[180] = chany_bottom_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[182];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[183];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[184] = chany_bottom_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[186];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[187];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[188] = chany_bottom_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[189] = chany_bottom_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[190] = chany_bottom_in[190];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[191] = chany_bottom_in[191];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[192] = chany_bottom_in[192];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[193] = chany_bottom_in[193];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[194] = chany_bottom_in[194];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[195] = chany_bottom_in[195];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[196] = chany_bottom_in[196];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[197] = chany_bottom_in[197];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[198] = chany_bottom_in[198];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[199] = chany_bottom_in[199];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[200] = chany_bottom_in[200];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[201] = chany_bottom_in[201];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[202] = chany_bottom_in[202];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[203] = chany_bottom_in[203];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[204] = chany_bottom_in[204];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[205] = chany_bottom_in[205];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[206] = chany_bottom_in[206];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[207] = chany_bottom_in[207];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[208] = chany_bottom_in[208];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[209] = chany_bottom_in[209];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[210] = chany_bottom_in[210];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[211] = chany_bottom_in[211];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[212] = chany_bottom_in[212];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[213] = chany_bottom_in[213];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[214] = chany_bottom_in[214];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[215] = chany_bottom_in[215];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[216] = chany_bottom_in[216];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[217] = chany_bottom_in[217];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[218] = chany_bottom_in[218];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[219] = chany_bottom_in[219];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[220] = chany_bottom_in[220];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[221] = chany_bottom_in[221];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[222] = chany_bottom_in[222];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[223] = chany_bottom_in[223];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[224] = chany_bottom_in[224];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[225] = chany_bottom_in[225];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[226] = chany_bottom_in[226];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[227] = chany_bottom_in[227];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[228] = chany_bottom_in[228];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[229] = chany_bottom_in[229];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[230] = chany_bottom_in[230];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[231] = chany_bottom_in[231];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[232] = chany_bottom_in[232];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[233] = chany_bottom_in[233];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[234] = chany_bottom_in[234];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[235] = chany_bottom_in[235];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[236] = chany_bottom_in[236];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[237] = chany_bottom_in[237];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[238] = chany_bottom_in[238];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[239] = chany_bottom_in[239];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[240] = chany_bottom_in[240];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[241] = chany_bottom_in[241];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[242] = chany_bottom_in[242];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[243] = chany_bottom_in[243];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[244] = chany_bottom_in[244];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[245] = chany_bottom_in[245];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[246] = chany_bottom_in[246];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[247] = chany_bottom_in[247];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[248] = chany_bottom_in[248];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[249] = chany_bottom_in[249];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[250] = chany_bottom_in[250];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[251] = chany_bottom_in[251];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[252] = chany_bottom_in[252];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[253] = chany_bottom_in[253];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[254] = chany_bottom_in[254];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[255] = chany_bottom_in[255];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[256] = chany_bottom_in[256];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[257] = chany_bottom_in[257];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[258] = chany_bottom_in[258];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[259] = chany_bottom_in[259];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[260] = chany_bottom_in[260];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[261] = chany_bottom_in[261];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[262] = chany_bottom_in[262];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[263] = chany_bottom_in[263];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[264] = chany_bottom_in[264];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[265] = chany_bottom_in[265];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[266] = chany_bottom_in[266];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[267] = chany_bottom_in[267];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[268] = chany_bottom_in[268];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[269] = chany_bottom_in[269];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[270] = chany_bottom_in[270];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[271] = chany_bottom_in[271];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[272] = chany_bottom_in[272];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[273] = chany_bottom_in[273];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[274] = chany_bottom_in[274];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[275] = chany_bottom_in[275];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[276] = chany_bottom_in[276];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[277] = chany_bottom_in[277];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[278] = chany_bottom_in[278];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[279] = chany_bottom_in[279];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[280] = chany_bottom_in[280];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[281] = chany_bottom_in[281];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[282] = chany_bottom_in[282];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[283] = chany_bottom_in[283];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[284] = chany_bottom_in[284];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[285] = chany_bottom_in[285];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[286] = chany_bottom_in[286];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[287] = chany_bottom_in[287];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[288] = chany_bottom_in[288];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[289] = chany_bottom_in[289];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[290] = chany_bottom_in[290];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[291] = chany_bottom_in[291];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[292] = chany_bottom_in[292];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[293] = chany_bottom_in[293];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[294] = chany_bottom_in[294];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[295] = chany_bottom_in[295];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[0] = chany_top_in[0];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[1];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[2];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[3];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[4] = chany_top_in[4];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[5];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[6];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[7];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[8] = chany_top_in[8];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[9];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[10];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[11];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[12] = chany_top_in[12];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[13];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[14];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[15];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[16] = chany_top_in[16];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[17];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[18];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[19];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[20] = chany_top_in[20];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[21];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[22];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[23];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[24] = chany_top_in[24];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[25];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[26];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[27];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[28] = chany_top_in[28];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[29];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[30];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[31];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[32] = chany_top_in[32];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[33];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[34];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[35];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[36] = chany_top_in[36];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[37];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[38];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[39];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[40] = chany_top_in[40];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[41];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[42];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[43];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[44] = chany_top_in[44];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[45];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[46];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[47];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[48] = chany_top_in[48];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[49];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[50];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[51];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[52] = chany_top_in[52];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[53];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[54];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[55];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[56] = chany_top_in[56];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[57];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[58];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[59];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[60] = chany_top_in[60];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[61];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[62];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[63];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[64] = chany_top_in[64];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[65] = chany_top_in[65];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[66] = chany_top_in[66];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[67] = chany_top_in[67];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[68] = chany_top_in[68];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chany_top_in[69];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[70] = chany_top_in[70];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[71] = chany_top_in[71];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[72] = chany_top_in[72];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[73] = chany_top_in[73];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[74] = chany_top_in[74];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[75] = chany_top_in[75];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[76] = chany_top_in[76];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[77] = chany_top_in[77];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[78] = chany_top_in[78];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[79] = chany_top_in[79];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[80] = chany_top_in[80];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[81] = chany_top_in[81];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[82] = chany_top_in[82];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[83] = chany_top_in[83];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[84] = chany_top_in[84];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[85] = chany_top_in[85];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[86] = chany_top_in[86];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[87] = chany_top_in[87];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[88] = chany_top_in[88];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[89] = chany_top_in[89];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[90] = chany_top_in[90];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[91] = chany_top_in[91];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[92] = chany_top_in[92];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[93] = chany_top_in[93];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[94] = chany_top_in[94];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[95] = chany_top_in[95];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[96] = chany_top_in[96];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[97] = chany_top_in[97];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[98] = chany_top_in[98];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[99] = chany_top_in[99];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[100] = chany_top_in[100];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[101] = chany_top_in[101];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[102] = chany_top_in[102];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[103] = chany_top_in[103];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[104] = chany_top_in[104];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[105] = chany_top_in[105];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[106] = chany_top_in[106];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[107] = chany_top_in[107];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[108] = chany_top_in[108];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[109] = chany_top_in[109];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[110] = chany_top_in[110];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[111] = chany_top_in[111];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[112] = chany_top_in[112];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[113] = chany_top_in[113];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[114] = chany_top_in[114];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[115] = chany_top_in[115];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[116] = chany_top_in[116];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[117] = chany_top_in[117];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[118] = chany_top_in[118];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[119] = chany_top_in[119];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[120] = chany_top_in[120];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[121] = chany_top_in[121];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[122] = chany_top_in[122];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[123] = chany_top_in[123];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[124] = chany_top_in[124];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[125] = chany_top_in[125];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[126] = chany_top_in[126];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[127] = chany_top_in[127];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[128] = chany_top_in[128];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[129] = chany_top_in[129];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[130] = chany_top_in[130];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[131] = chany_top_in[131];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[132] = chany_top_in[132];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[133] = chany_top_in[133];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[134] = chany_top_in[134];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[135] = chany_top_in[135];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[136] = chany_top_in[136];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[137] = chany_top_in[137];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[138] = chany_top_in[138];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[139] = chany_top_in[139];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[140] = chany_top_in[140];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[141] = chany_top_in[141];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[142] = chany_top_in[142];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[143] = chany_top_in[143];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[144] = chany_top_in[144];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[145] = chany_top_in[145];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[146] = chany_top_in[146];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[147] = chany_top_in[147];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[148] = chany_top_in[148];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[149] = chany_top_in[149];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[150] = chany_top_in[150];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[151] = chany_top_in[151];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[152] = chany_top_in[152];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[153] = chany_top_in[153];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[154] = chany_top_in[154];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[155] = chany_top_in[155];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[156] = chany_top_in[156];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[157] = chany_top_in[157];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[158] = chany_top_in[158];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[159] = chany_top_in[159];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[160] = chany_top_in[160];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[161] = chany_top_in[161];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[162] = chany_top_in[162];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[163] = chany_top_in[163];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[164] = chany_top_in[164];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[165] = chany_top_in[165];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[166] = chany_top_in[166];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[167] = chany_top_in[167];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[168] = chany_top_in[168];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[169] = chany_top_in[169];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[170] = chany_top_in[170];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[171] = chany_top_in[171];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[172] = chany_top_in[172];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[173] = chany_top_in[173];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[174] = chany_top_in[174];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[175] = chany_top_in[175];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[176] = chany_top_in[176];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[177] = chany_top_in[177];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[178] = chany_top_in[178];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[179] = chany_top_in[179];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[180] = chany_top_in[180];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[181] = chany_top_in[181];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[182] = chany_top_in[182];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[183] = chany_top_in[183];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[184] = chany_top_in[184];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[185] = chany_top_in[185];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[186] = chany_top_in[186];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[187] = chany_top_in[187];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[188] = chany_top_in[188];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[189] = chany_top_in[189];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[190] = chany_top_in[190];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[191] = chany_top_in[191];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[192] = chany_top_in[192];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[193] = chany_top_in[193];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[194] = chany_top_in[194];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[195] = chany_top_in[195];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[196] = chany_top_in[196];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[197] = chany_top_in[197];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[198] = chany_top_in[198];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[199] = chany_top_in[199];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[200] = chany_top_in[200];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[201] = chany_top_in[201];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[202] = chany_top_in[202];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[203] = chany_top_in[203];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[204] = chany_top_in[204];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[205] = chany_top_in[205];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[206] = chany_top_in[206];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[207] = chany_top_in[207];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[208] = chany_top_in[208];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[209] = chany_top_in[209];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[210] = chany_top_in[210];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[211] = chany_top_in[211];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[212] = chany_top_in[212];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[213] = chany_top_in[213];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[214] = chany_top_in[214];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[215] = chany_top_in[215];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[216] = chany_top_in[216];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[217] = chany_top_in[217];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[218] = chany_top_in[218];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[219] = chany_top_in[219];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[220] = chany_top_in[220];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[221] = chany_top_in[221];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[222] = chany_top_in[222];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[223] = chany_top_in[223];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[224] = chany_top_in[224];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[225] = chany_top_in[225];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[226] = chany_top_in[226];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[227] = chany_top_in[227];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[228] = chany_top_in[228];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[229] = chany_top_in[229];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[230] = chany_top_in[230];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[231] = chany_top_in[231];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[232] = chany_top_in[232];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[233] = chany_top_in[233];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[234] = chany_top_in[234];
// ----- Local connection due to Wire 531 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[235] = chany_top_in[235];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[236] = chany_top_in[236];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[237] = chany_top_in[237];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[238] = chany_top_in[238];
// ----- Local connection due to Wire 535 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[239] = chany_top_in[239];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[240] = chany_top_in[240];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[241] = chany_top_in[241];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[242] = chany_top_in[242];
// ----- Local connection due to Wire 539 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[243] = chany_top_in[243];
// ----- Local connection due to Wire 540 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[244] = chany_top_in[244];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[245] = chany_top_in[245];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[246] = chany_top_in[246];
// ----- Local connection due to Wire 543 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[247] = chany_top_in[247];
// ----- Local connection due to Wire 544 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[248] = chany_top_in[248];
// ----- Local connection due to Wire 545 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[249] = chany_top_in[249];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[250] = chany_top_in[250];
// ----- Local connection due to Wire 547 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[251] = chany_top_in[251];
// ----- Local connection due to Wire 548 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[252] = chany_top_in[252];
// ----- Local connection due to Wire 549 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[253] = chany_top_in[253];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[254] = chany_top_in[254];
// ----- Local connection due to Wire 551 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[255] = chany_top_in[255];
// ----- Local connection due to Wire 552 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[256] = chany_top_in[256];
// ----- Local connection due to Wire 553 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[257] = chany_top_in[257];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[258] = chany_top_in[258];
// ----- Local connection due to Wire 555 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[259] = chany_top_in[259];
// ----- Local connection due to Wire 556 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[260] = chany_top_in[260];
// ----- Local connection due to Wire 557 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[261] = chany_top_in[261];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[262] = chany_top_in[262];
// ----- Local connection due to Wire 559 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[263] = chany_top_in[263];
// ----- Local connection due to Wire 560 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[264] = chany_top_in[264];
// ----- Local connection due to Wire 561 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[265] = chany_top_in[265];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[266] = chany_top_in[266];
// ----- Local connection due to Wire 563 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[267] = chany_top_in[267];
// ----- Local connection due to Wire 564 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[268] = chany_top_in[268];
// ----- Local connection due to Wire 565 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[269] = chany_top_in[269];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[270] = chany_top_in[270];
// ----- Local connection due to Wire 567 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[271] = chany_top_in[271];
// ----- Local connection due to Wire 568 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[272] = chany_top_in[272];
// ----- Local connection due to Wire 569 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[273] = chany_top_in[273];
// ----- Local connection due to Wire 570 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[274] = chany_top_in[274];
// ----- Local connection due to Wire 571 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[275] = chany_top_in[275];
// ----- Local connection due to Wire 572 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[276] = chany_top_in[276];
// ----- Local connection due to Wire 573 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[277] = chany_top_in[277];
// ----- Local connection due to Wire 574 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[278] = chany_top_in[278];
// ----- Local connection due to Wire 575 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[279] = chany_top_in[279];
// ----- Local connection due to Wire 576 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[280] = chany_top_in[280];
// ----- Local connection due to Wire 577 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[281] = chany_top_in[281];
// ----- Local connection due to Wire 578 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[282] = chany_top_in[282];
// ----- Local connection due to Wire 579 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[283] = chany_top_in[283];
// ----- Local connection due to Wire 580 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[284] = chany_top_in[284];
// ----- Local connection due to Wire 581 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[285] = chany_top_in[285];
// ----- Local connection due to Wire 582 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[286] = chany_top_in[286];
// ----- Local connection due to Wire 583 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[287] = chany_top_in[287];
// ----- Local connection due to Wire 584 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[288] = chany_top_in[288];
// ----- Local connection due to Wire 585 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[289] = chany_top_in[289];
// ----- Local connection due to Wire 586 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[290] = chany_top_in[290];
// ----- Local connection due to Wire 587 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[291] = chany_top_in[291];
// ----- Local connection due to Wire 588 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[292] = chany_top_in[292];
// ----- Local connection due to Wire 589 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[293] = chany_top_in[293];
// ----- Local connection due to Wire 590 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[294] = chany_top_in[294];
// ----- Local connection due to Wire 591 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[295] = chany_top_in[295];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size100 mux_left_ipin_0 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_0_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_0_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_0_));

	mux_tree_tapbuf_size100 mux_left_ipin_1 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_1_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_1_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_1_));

	mux_tree_tapbuf_size100 mux_left_ipin_2 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_2_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_2_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_2_));

	mux_tree_tapbuf_size100 mux_left_ipin_3 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_3_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_3_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_3_));

	mux_tree_tapbuf_size100 mux_left_ipin_4 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_4_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_4_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_4_));

	mux_tree_tapbuf_size100 mux_left_ipin_5 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_5_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_5_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_5_));

	mux_tree_tapbuf_size100 mux_left_ipin_6 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_6_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_6_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_6_));

	mux_tree_tapbuf_size100 mux_left_ipin_7 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_7_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_7_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_7_));

	mux_tree_tapbuf_size100 mux_left_ipin_8 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_8_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_8_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_8_));

	mux_tree_tapbuf_size100 mux_left_ipin_9 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_9_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_9_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_9_));

	mux_tree_tapbuf_size100 mux_left_ipin_10 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_10_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_10_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_10_));

	mux_tree_tapbuf_size100 mux_left_ipin_11 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_11_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_11_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_11_));

	mux_tree_tapbuf_size100 mux_left_ipin_12 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_12_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_12_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_12_));

	mux_tree_tapbuf_size100 mux_left_ipin_13 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_13_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_13_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_13_));

	mux_tree_tapbuf_size100 mux_left_ipin_14 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_14_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_14_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_14_));

	mux_tree_tapbuf_size100 mux_left_ipin_15 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_15_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_15_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_15_));

	mux_tree_tapbuf_size100 mux_left_ipin_16 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_16_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_16_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_16_));

	mux_tree_tapbuf_size100 mux_left_ipin_17 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_17_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_17_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_17_));

	mux_tree_tapbuf_size100 mux_left_ipin_18 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_18_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_18_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_18_));

	mux_tree_tapbuf_size100 mux_left_ipin_19 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_19_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_19_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_19_));

	mux_tree_tapbuf_size100 mux_left_ipin_20 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_20_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_20_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_20_));

	mux_tree_tapbuf_size100 mux_left_ipin_21 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_21_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_21_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_21_));

	mux_tree_tapbuf_size100 mux_left_ipin_22 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_22_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_22_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_22_));

	mux_tree_tapbuf_size100 mux_left_ipin_23 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_23_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_23_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_23_));

	mux_tree_tapbuf_size100 mux_left_ipin_24 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_24_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_24_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_24_));

	mux_tree_tapbuf_size100 mux_left_ipin_25 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_25_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_25_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_25_));

	mux_tree_tapbuf_size100 mux_left_ipin_26 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_26_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_26_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_26_));

	mux_tree_tapbuf_size100 mux_left_ipin_27 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_27_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_27_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_27_));

	mux_tree_tapbuf_size100 mux_left_ipin_28 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_28_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_28_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_28_));

	mux_tree_tapbuf_size100 mux_left_ipin_29 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_29_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_29_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_29_));

	mux_tree_tapbuf_size100 mux_left_ipin_30 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_30_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_30_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_30_));

	mux_tree_tapbuf_size100 mux_left_ipin_31 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_31_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_31_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_31_));

	mux_tree_tapbuf_size100 mux_left_ipin_32 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_32_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_32_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_32_));

	mux_tree_tapbuf_size100 mux_left_ipin_33 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_33_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_33_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_33_));

	mux_tree_tapbuf_size100 mux_left_ipin_34 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_34_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_34_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_34_));

	mux_tree_tapbuf_size100 mux_left_ipin_35 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_35_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_35_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_35_));

	mux_tree_tapbuf_size100 mux_left_ipin_36 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_36_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_36_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_36_));

	mux_tree_tapbuf_size100 mux_left_ipin_37 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_37_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_37_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_37_));

	mux_tree_tapbuf_size100 mux_left_ipin_38 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_38_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_38_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_38_));

	mux_tree_tapbuf_size100 mux_left_ipin_39 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_39_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_39_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_39_));

	mux_tree_tapbuf_size100 mux_left_ipin_40 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_40_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_40_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_40_));

	mux_tree_tapbuf_size100 mux_left_ipin_41 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_41_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_41_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_41_));

	mux_tree_tapbuf_size100 mux_left_ipin_42 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_42_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_42_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_42_));

	mux_tree_tapbuf_size100 mux_left_ipin_43 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_43_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_43_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_43_));

	mux_tree_tapbuf_size100 mux_left_ipin_44 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_44_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_44_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_44_));

	mux_tree_tapbuf_size100 mux_left_ipin_45 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_45_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_45_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_45_));

	mux_tree_tapbuf_size100 mux_left_ipin_46 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_46_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_46_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_46_));

	mux_tree_tapbuf_size100 mux_left_ipin_47 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_47_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_47_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_47_));

	mux_tree_tapbuf_size100 mux_left_ipin_48 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_48_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_48_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_48_));

	mux_tree_tapbuf_size100 mux_left_ipin_49 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_49_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_49_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_49_));

	mux_tree_tapbuf_size100 mux_left_ipin_50 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_50_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_50_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_50_));

	mux_tree_tapbuf_size100 mux_left_ipin_51 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_51_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_51_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_51_));

	mux_tree_tapbuf_size100 mux_left_ipin_52 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_52_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_52_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_52_));

	mux_tree_tapbuf_size100 mux_left_ipin_53 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_53_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_53_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_53_));

	mux_tree_tapbuf_size100 mux_left_ipin_54 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_54_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_54_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_54_));

	mux_tree_tapbuf_size100 mux_left_ipin_55 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_55_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_55_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_55_));

	mux_tree_tapbuf_size100 mux_left_ipin_56 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_56_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_56_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_56_));

	mux_tree_tapbuf_size100 mux_left_ipin_57 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_57_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_57_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_57_));

	mux_tree_tapbuf_size100 mux_left_ipin_58 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_58_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_58_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_58_));

	mux_tree_tapbuf_size100 mux_left_ipin_59 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_59_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_59_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_59_));

	mux_tree_tapbuf_size100 mux_left_ipin_60 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_60_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_60_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_60_));

	mux_tree_tapbuf_size100 mux_left_ipin_61 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_61_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_61_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_61_));

	mux_tree_tapbuf_size100 mux_left_ipin_62 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_62_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_62_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_62_));

	mux_tree_tapbuf_size100 mux_left_ipin_63 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_63_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_63_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_63_));

	mux_tree_tapbuf_size100 mux_left_ipin_64 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_64_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_64_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_64_));

	mux_tree_tapbuf_size100 mux_left_ipin_65 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_65_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_65_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_65_));

	mux_tree_tapbuf_size100 mux_left_ipin_66 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_66_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_66_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_66_));

	mux_tree_tapbuf_size100 mux_left_ipin_67 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_67_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_67_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_67_));

	mux_tree_tapbuf_size100 mux_left_ipin_68 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_68_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_68_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_68_));

	mux_tree_tapbuf_size100 mux_left_ipin_69 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_69_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_69_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_3_69_));

	mux_tree_tapbuf_size100 mux_left_ipin_70 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_70_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_70_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_0_));

	mux_tree_tapbuf_size100 mux_left_ipin_71 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_71_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_71_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_1_));

	mux_tree_tapbuf_size100 mux_left_ipin_72 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_72_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_72_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_2_));

	mux_tree_tapbuf_size100 mux_left_ipin_73 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187], chany_bottom_in[193], chany_top_in[193], chany_bottom_in[199], chany_top_in[199], chany_bottom_in[205], chany_top_in[205], chany_bottom_in[211], chany_top_in[211], chany_bottom_in[217], chany_top_in[217], chany_bottom_in[223], chany_top_in[223], chany_bottom_in[229], chany_top_in[229], chany_bottom_in[235], chany_top_in[235], chany_bottom_in[241], chany_top_in[241], chany_bottom_in[247], chany_top_in[247], chany_bottom_in[253], chany_top_in[253], chany_bottom_in[259], chany_top_in[259], chany_bottom_in[265], chany_top_in[265], chany_bottom_in[271], chany_top_in[271], chany_bottom_in[277], chany_top_in[277], chany_bottom_in[283], chany_top_in[283], chany_bottom_in[289], chany_top_in[289], chany_bottom_in[295], chany_top_in[295]}),
		.sram(mux_tree_tapbuf_size100_73_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_73_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_0_));

	mux_tree_tapbuf_size100 mux_left_ipin_74 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188], chany_bottom_in[194], chany_top_in[194], chany_bottom_in[200], chany_top_in[200], chany_bottom_in[206], chany_top_in[206], chany_bottom_in[212], chany_top_in[212], chany_bottom_in[218], chany_top_in[218], chany_bottom_in[224], chany_top_in[224], chany_bottom_in[230], chany_top_in[230], chany_bottom_in[236], chany_top_in[236], chany_bottom_in[242], chany_top_in[242], chany_bottom_in[248], chany_top_in[248], chany_bottom_in[254], chany_top_in[254], chany_bottom_in[260], chany_top_in[260], chany_bottom_in[266], chany_top_in[266], chany_bottom_in[272], chany_top_in[272], chany_bottom_in[278], chany_top_in[278], chany_bottom_in[284], chany_top_in[284], chany_bottom_in[290], chany_top_in[290]}),
		.sram(mux_tree_tapbuf_size100_74_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_74_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_1_));

	mux_tree_tapbuf_size100 mux_left_ipin_75 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183], chany_bottom_in[189], chany_top_in[189], chany_bottom_in[195], chany_top_in[195], chany_bottom_in[201], chany_top_in[201], chany_bottom_in[207], chany_top_in[207], chany_bottom_in[213], chany_top_in[213], chany_bottom_in[219], chany_top_in[219], chany_bottom_in[225], chany_top_in[225], chany_bottom_in[231], chany_top_in[231], chany_bottom_in[237], chany_top_in[237], chany_bottom_in[243], chany_top_in[243], chany_bottom_in[249], chany_top_in[249], chany_bottom_in[255], chany_top_in[255], chany_bottom_in[261], chany_top_in[261], chany_bottom_in[267], chany_top_in[267], chany_bottom_in[273], chany_top_in[273], chany_bottom_in[279], chany_top_in[279], chany_bottom_in[285], chany_top_in[285], chany_bottom_in[291], chany_top_in[291]}),
		.sram(mux_tree_tapbuf_size100_75_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_75_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_2_));

	mux_tree_tapbuf_size100 mux_right_ipin_0 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184], chany_bottom_in[190], chany_top_in[190], chany_bottom_in[196], chany_top_in[196], chany_bottom_in[202], chany_top_in[202], chany_bottom_in[208], chany_top_in[208], chany_bottom_in[214], chany_top_in[214], chany_bottom_in[220], chany_top_in[220], chany_bottom_in[226], chany_top_in[226], chany_bottom_in[232], chany_top_in[232], chany_bottom_in[238], chany_top_in[238], chany_bottom_in[244], chany_top_in[244], chany_bottom_in[250], chany_top_in[250], chany_bottom_in[256], chany_top_in[256], chany_bottom_in[262], chany_top_in[262], chany_bottom_in[268], chany_top_in[268], chany_bottom_in[274], chany_top_in[274], chany_bottom_in[280], chany_top_in[280], chany_bottom_in[286], chany_top_in[286], chany_bottom_in[292], chany_top_in[292]}),
		.sram(mux_tree_tapbuf_size100_76_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_76_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_I_1_));

	mux_tree_tapbuf_size100 mux_right_ipin_1 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185], chany_bottom_in[191], chany_top_in[191], chany_bottom_in[197], chany_top_in[197], chany_bottom_in[203], chany_top_in[203], chany_bottom_in[209], chany_top_in[209], chany_bottom_in[215], chany_top_in[215], chany_bottom_in[221], chany_top_in[221], chany_bottom_in[227], chany_top_in[227], chany_bottom_in[233], chany_top_in[233], chany_bottom_in[239], chany_top_in[239], chany_bottom_in[245], chany_top_in[245], chany_bottom_in[251], chany_top_in[251], chany_bottom_in[257], chany_top_in[257], chany_bottom_in[263], chany_top_in[263], chany_bottom_in[269], chany_top_in[269], chany_bottom_in[275], chany_top_in[275], chany_bottom_in[281], chany_top_in[281], chany_bottom_in[287], chany_top_in[287], chany_bottom_in[293], chany_top_in[293]}),
		.sram(mux_tree_tapbuf_size100_77_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_77_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_I_5_));

	mux_tree_tapbuf_size100 mux_right_ipin_2 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186], chany_bottom_in[192], chany_top_in[192], chany_bottom_in[198], chany_top_in[198], chany_bottom_in[204], chany_top_in[204], chany_bottom_in[210], chany_top_in[210], chany_bottom_in[216], chany_top_in[216], chany_bottom_in[222], chany_top_in[222], chany_bottom_in[228], chany_top_in[228], chany_bottom_in[234], chany_top_in[234], chany_bottom_in[240], chany_top_in[240], chany_bottom_in[246], chany_top_in[246], chany_bottom_in[252], chany_top_in[252], chany_bottom_in[258], chany_top_in[258], chany_bottom_in[264], chany_top_in[264], chany_bottom_in[270], chany_top_in[270], chany_bottom_in[276], chany_top_in[276], chany_bottom_in[282], chany_top_in[282], chany_bottom_in[288], chany_top_in[288], chany_bottom_in[294], chany_top_in[294]}),
		.sram(mux_tree_tapbuf_size100_78_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size100_78_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_I_9_));

	mux_tree_tapbuf_size100_mem mem_left_ipin_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size100_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_0_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_0_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_1_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_1_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_2_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_2_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_3_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_3_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_4_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_4_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_5_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_5_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_6_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_6_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_7_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_7_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_8_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_8_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_9_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_9_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_10_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_10_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_11_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_11_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_12_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_12_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_13_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_13_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_14_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_14_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_15_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_15_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_16_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_16_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_17_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_17_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_18_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_18_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_19_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_19_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_20_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_20_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_21_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_21_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_22_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_22_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_23_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_23_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_24_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_24_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_25_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_25_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_26_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_26_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_27_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_27_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_28_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_28_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_29_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_29_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_30_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_30_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_31_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_31_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_32_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_32_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_33_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_33_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_34_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_34_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_35_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_35_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_36_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_36_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_37_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_37_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_38_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_38_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_39_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_39_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_40_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_40_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_41_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_41_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_42_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_42_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_43_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_43_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_44_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_44_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_45_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_45_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_46_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_46_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_47_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_47_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_48_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_48_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_49_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_49_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_50_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_50_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_51_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_51_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_52_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_52_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_53_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_53_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_54_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_54_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_55_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_55_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_56_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_56_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_57_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_57_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_58_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_58_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_59_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_59_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_60_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_60_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_61_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_61_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_62_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_62_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_63_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_63_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_64_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_64_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_65_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_65_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_66_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_66_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_67_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_67_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_68_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_68_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_69_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_69_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_70_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_70_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_71_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_71_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_72_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_72_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_73_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_73_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_74_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_74_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_left_ipin_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_75_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_75_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_right_ipin_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_76_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_76_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_right_ipin_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size100_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_77_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_77_sram_inv[0:6]));

	mux_tree_tapbuf_size100_mem mem_right_ipin_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size100_mem_77_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size100_78_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size100_78_sram_inv[0:6]));

endmodule
// ----- END Verilog module for cby_5__6_ -----

//----- Default net type -----
`default_nettype wire




